//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Tzu-Yun Huang
//	 Editor		: Ting-Yu Chang
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_DRAM.v
//   Module Name : pseudo_DRAM
//   Release version : v3.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module pseudo_DRAM
`protected
(?c^L3AR4g,QTc?f,H##TN;LK]N:.H]D2UQ]g&9Kb(cU(J/,PU#R-)_X9=?O&5da
+2\B^RLf8fS_gXV8/LN-_>@Bb_^6;2YZ=;WP=A6^BJ>d]23f9d^QNF=>fY2C;JC[
[V_NK5dV<&R6JGAI2ZIHMQEYWF.W17E&1>(EBF9(K=FB_S^[^OGCXF>>8&G2G@E0
dP88;8QLJad)CdaE9:BOREd8Z<J_&g<P0(7M,7/E60?-,<PCY[LM5.[cDJbI4TOW
W+eBM<RE[R]=I5c34:@X]AbQd1+(c3H^a8Q6cc)-7QR4^(?;HAJg06T;BE,ZWeBP
#>cBWVF;FQ##TEK+)_f(80O2_B0/bJOg,K5&M04e)J_#V5L]9/+)W^[e^1VdVPgR
<@-6^4(J54]M0[>-MV&dG0/5N@;ED9JH_d[AH.2<=6H<ET^M#D86-@<U3)#-A=2c
eEZ_-[4+T2+R(B40W?6UAaDM</c)K3H0AT]YJ[641FJN?eY=Ad>[.7S;24,&2gE]
Db&UVWSC<cB^(Lg(@V&LEV2V=KAU^CGS2YH#V+BOX8H&;FUa&REdZJ,08cR0U=V1
WXDF0/L/#C.J=L;C4K>1-,Q;RHSTf[]>PSa2BG]<OGW9+Q7-<WFKI&>N.NGWNY&M
YC\9Q+a6.c\U1@Ve0Z(I[ESa;b)Gb5gZG/RI^[Q<NO)E]DB5bgND>b>^HYNC_QB&
QZF+7FH8/4&3M^Z5,1\&Z])(/I0#.9[:+S9I6QFGQ^M\Q:4TP3(M9V5B@/ZV,6\5
PUfOL)?3dKMZ<cZU8g<)T^2B4)LDSJ&NaRNKW=H1e\\2F8EL:]eFF;WSSdg&:5?f
Z4DCF[[@9X&BC](g.fH7<_-\E\bYe9:1]K8Y-3-G@XBCD&>/5(Y0=Ug8Y5B=1?Qc
42JJD)NO&_A^SVHe<+#)08?Q-FZ#,aBZfY>+^_NU<_ef?ROf\=?[Bg,5UIbQ8.Z?
#T_+-M4BFQ?MFV.3,2HfVS+YX1KA\9EMa/[5AP5J8Z&,cYKgCF#V9&E-3_V_VG0.
I&#95?^gQ1IA6dFSZ]Ydg1RMId0+9=;bU?]c\Y8Q]U5>.5bdPRM(cOH^I#[XD)[U
T,,5bS#PEa2:GL>3dg-.G+.NN[EeI6c[J^c)JFYA;6DGV1Ya:L#e37A_\?(YW8J:
Jc7Vc1J5-ES#a.aMDUd#GZG&E>M9R#]VcZ][d7GP2Y-;O[5=;IJ7=@?A+\\Zbg)O
Ag&VT84aQ^T+_D?+HLJ+TQW0O?ggeTfG(.:+ALgK]aMV2Ma+=@B,IHNYI/]XUZ:G
?XL6K;C:V@LL>a,=TW[SDV,e19A,4^GaZ>WWc8A?gL\]9PRS/;+T;F-;cIAF&Y(O
D[bJc7;K0Mb3,6Db#8((BOXG?I4D/6TV@H@9d\3KG]Q)@9HT:7G8-4aOIX&VI=FP
7EeCgg];^bD8B.S2V3U8=EUCYDZZ_U\7,:&_cc(EMROSY;(U#6N;QQW,W:8.e.M=
\YfeZgQH7([Z/KB\724-@VffK(M8&<g@[8NRWN0DQF=T,:7K_39@(FT:#:F8\@/U
>H_2\.31B9fIGH:VK]KJW53\,4,^06AUE+AeSJBO9c9&23@3(EDM#fUf0:GHd5R9
RS0.PYAFH:M4_63^bgK:Cg34\f<#\]M9X7Z.1:GC@3ga^2Xe^BgT6b<R-3a)?0AE
V<J5,HZ+ODT>e?^<)-@C?:]c4IC@b]O-Nf.DN,5(WO-5)N_0bSF^.:G=TEXINd;g
40R6?#G+=(H/aeBXVAS3HL2<)aY[GP8BSGE88GKL^]BEZL;G&T?_/[DP/)GQ:Q;F
2PFa5RA1NQN2+)EGPB8T\,QJ,MBGP)BM9SN_OT]W0:]dA5+O3UH0(0GZD=ScYO]_
&7L>dWHf8R&&RSbT_MYEL/^HXRX\9Y^9UB6._J.-)Td/XJ@b4Zc5&3X9?B94K9Ud
OI4#G1b@U-S#<G#^2D?0R4T6HPY()a0P0P?^Z>;?YfCVRHL?[KHQ[:.-O#Z-a=Z@
eX/:=Ya34G>U1YgYR1.<(>;M&\FFA<9+-6AU/-4I@L13NR46\O+Rf)T4egIg_X3g
d/Jc:;D2>:GK9GFU:f/(YY:&-Z]PSH8_N:&SO29Z^]80Z^0H(H2=_@ILA&#4.Lc9
6TE[g(U^2?&d@Z)THH>I,3A;6a;LMWb8K0;4@-dVgM:=Z1Q2@<3?-GA^DG8a3B2\
Zf)eJF\e3b[EZ:be4]VD]=868S0;+d6,I,Z1MQe&6e0KUQ#^P?47d_(RP-c)GT5d
=UXPGGYL1:JK;bHY??Y/d?LZ8c#Y^=X>_\5Td4W_&VEG=<O7.U3(Wg2ZXff_#\D+
dbI(bd.XKe2Z,R/4gR[WJGN+\Z>)1dU.JI+dO;V01P(=cF.\#X?VPgFSQ)F/XTeV
gM7VR\SNA=b9eI_QV7,TFZ@YT\NHGaM1HE=MG;;0<0,O1D<EE.\^0C)]+<76)Mga
GG_/d]7Vd-a6>+I0P^NRL64Kf9L8+3QfWO#fT)),\0,9JM+eB&1f\EgTU8E9.)b4
-ENP7MO(<^FT:F^gCJf5E1IZN_g6Fc;?KP<\0B#3Q^-MNCMeD7&X3V2JH:_K>dS(
0:cWWTKXe>2\DV4;&QYfEOJK(YGX\[[C/5L>LZWZ4^:@:1d[2UL&YC63)SNg.:A(
cF0S/5Q(16dNQ_a2Ua;(D898#]3GC[=@R^^GfB3V=)J#<3\GL9M/-EH=b=IMag9Q
dAX1,,c,M=2(XeJG>?-XZR\5#XUaU5WH6NefWN<e(eM<6^c60b\-Z=-_Q7<JgA/f
6#WZBHB>DCY@6c\=gfd3QPRdV.d=VH#[C5OIa6/\0aW=3>T:X/42=6UPHS)W@P_G
Db.:#e+DX:YPHa;FQ;\eM/eCUV-a^XC=#P5_E:.PcGS\P83UTM#-&-\B-8NT&QTR
&0e#6S4)B2-[(3B=X_GUS1&9@2_ZJ]M-]P9FY/OWT>_)9YYN]ReCMf8L&<P2BV7d
K0LPTVX+ANaFR6T<6N5:Q#E+VD&K;BS,BXV8T[fc.4I^\/;B6NUH.0[=LRY?:6L/
OK5cb?>)KFQ,MX+]2UJQ:-0cV=8]a=IOJV[.(@,O(-:<?.F5K4D>/bZ];8_M;Y^B
:RE]Qc&.R-9-cbXe.:FfLKOFROV3A@L_4J)H440:dBe[63&D1^RLGZKd^Y=:AZ;(
cW@N>8eg,GKe:\=JVCbOGdgU+=>\6T2_RR\7UY:C&<0-cL<7gddS;A;1\2_5M9e,
e)L]19;Fg(?CL+FRTbEZU6-X>[4eG@8S.QG1\L\7W:5GJ/\JFX+B2d5b9_DM5,Ua
Y[5HPB<LIR8.RbQWN72RB&:adG.SP2#\4]2+#g+:ZGbgD&?V12<P^VdOEg_MH4[L
#EEMO^X1XfJ><I5#5GF7B&<:34^AgCDYEKFIA_FOTC0GBCLQM@cKX=Q;dXI)Q>\f
WB_(gQ(,R<D7TM5OT07WVO21=_bI:P\:ed=Y;fM&X]e4+,<&Xf)C4.HGag8O0LLZ
U9]DPcDTAXBW?g\@,)2&#VP]OQS@_S]VK2\R<R/WGVMEYPJXB3^Ob50DLg.L^M-4
^.^[BBaaL,DS[R@+^.EZIe2e^;T?6ZMf?Q\4:G:,7-\PW;;Cg-g]U_0\c1d.5-3Q
Y@LCP7f7@g^VCVZZ.b,d>Bd\,L_bO)SdaXKA9EWS31gFO=<W,[Q5c>R.?@HJ\Q=c
K;.&DTZ;>@6+Ba#ZU8#J4Wce^Ve3@VD<-)2\2gG2g9:(T8YPCZD2N<3bXZ_L7W2.
KgZA)fcA4d7N9.5D[J2fEYM58@caRV(_2BBRP2G1_7CD6U7P+C?8)YN8GdH4=1UO
?60Z&<d+(3ZDLJ=N>P[1Eaa4#-9OU=OaQR8LJ.ZWE?Y?U@09>JIJN84M)K7J5CY>
MgBG;02A@6BKfbDd>4L,753NHD9Md(d_4HM7a^5f7B21_ZXGSQ^J:;,_Y;#=<_8G
H/IU7+YK0909WD>,a-M^<K^Q16TQ??3GE8_QE,2ZZ-V8ISEWe[\dc,f7B3A1KNH?
:HO]EFgfG3/V@@=bg,4IJV,6Q^S.^:&<14AC)\N&N<<H83dLSdD@I=.a+7+W(RQQ
Z]BXbEGB1Zg\))2E]0^XQCKP13=XdDYY7I;cQ5XURA:4=-QV@e9+6,K_US;-^+F,
5X+^gJM&DUMab;P+_(]IBO@=@Y6g=R#fUVG\D]DWgbG30\2&N+D:;(CSL\X-HdHL
G6ZGgb]8U<8)5bg;N<9=LP789\0Z5MX_E]Zb[&@CTTWIC^+C&JBJ+1LIC@M8_3[,
K66OV_fLNa\7(]C6c^)\]1Y/#2D<PW36(C(CVA]JLJcV+Z2Mb1+4g]JILE[XWEVD
AbX_14&_+@D(6CKD4)O6:/27(;7O=<Z3AKT-TF0P5?TNT.<gWeC8\/F#?]VL:-S-
CgR\UP)e+T/2CR=O(25:Kc2<gPKc&gSA6?;S(bb40E]N16L,f2R#)OY0LNFR&Z(Z
@0A9[cD66cKYZ)IUdaLS3=TEDV,/A?XTQ+_K:4DCP@e1,&__W^?C^U/2T,Gd=Gg0
+d+f-YbgR-2H[Sbb(W:#O,-UO.V1.FId_7gWI[gT+O(M13E\:VAY8A9d<?a1RT;X
>5B1g?Q6-3@,)FG2SDQ@JN(F7VRT788K5-SLC4#c2GNJ_Z/X[8BF0R\KbOHb/_FU
^SNQ=CODZY^>58bK?Db62Ha-3?U)V+S&&9dS/KYI[BMQ9HZ)9=6FX3_M<_KDGR&#
d:<00JDV+CP>V7F1T06/SJ\.[Hed1CJ1#;/f2ee5PT0+O5ZUO0IR(fL)]-(;+?dI
KGLKST.2;5T>S/2f-56<.NRA\bG=#T,+N3,VOJB.-O;6b<R39?YGNSRFFa1HcNV;
F?].UGHA]1WX-fPdZA4P&X/UGE.0=QKKdJ#4+#/_OP6,HIdJ/FKe//Yd=OV:=6:M
(c437H207MX5J,gAMV#.7+MOTd=d\^[ZeA)>Q,P&Q\]O@S<5U7_0<L)_8)@/d@#<
CbCbYC;U1V3-GCOH\O>,>;B&T#CNd7?=CN4U_P9?=5JZ8d\)d#FA#;?)8g&eZ_V.
VP/fD^_JH=50d9I8.RNHRS(7#_7DGZNCNLJWgNeB<MG[Z7\.E+b56Lf&>,f2_YfI
5WAeHP^2+?YcC/eLS9N,LKX\eXf.88g@AM<1K8LM4Q=;=ac_+Ec^T=Q,9B)QRaS3
Y:6Rc57WA)ZOK;&V)F60\Sa.^#^AceOQ\b._Y_&fL(O7>;,.&]M-Q,&Kf,Z13.?_
0,#,[0[QG]9M)RKEa(EI:cRgF#Q7]L<Q=C\[(#YV&A+>18Q__]7@A]/PL&K(LDU5
IMBFg-07UN,][aZ+)@MI=^[A(&eE46>N@G&XC(<RK),(Q5cNU2-G3I76&^Y8Z5^(
1=1+\)?aWP6)JY\&=MJ<\7c6f2H1(];d74&\).c]RK63GIC3U#8e,fY@?g:?)<a>
>9N6/.377PW:+d>K+09O<ZHOZ@><C^+5]:F7^e3EO.[GD9W1ES-afE1;)?5/H7af
@_7G:F\K>U^Tf0gII^(AecG?U?CFOAZ5LU,J@=.9P[6d<J_NC=&bI+>W/AaZ36BU
76H^7G?3GL@7_C6QOM5IZ?X.KHdK@C4,YgU:5DO8bI]Qe6?T93/5P<9\^bH5Z.+>
&-@XTN3<>-V=1DLLM]A\97U0ZDS2QD-83bbaM4(+^SYV7(A.6<O.Gb[O@AFQL]XL
/L2;bQZ]E]92I]7>e#3_GCZM3J(KGRGV0((BW.<:&\;g1P70OO+@^W&cFJV.P+-:
RL>f^eQ4N^fEI1/aF6HI=;_?Y3I4@N^0]Nf7@eU&(T>a)97;d1-4eODE@_FDT.L6
@f9G)&>X58PdJ#&:Q<3QZb<<I:ge0-(CTc)I:4.)=.a3FEZ-V^SIf?ZZ72^BGS7Q
M)AaCJIeM2c5Q?KN&CPFT=8^fdY7H1XVPYWX5cH)(O(5NPGJ:J1Ma40g(Y#5/T,O
/5d7^^8G[W4T;&B\c#^]5Y,PSH-H#eNN8dG7>:W_/_a9+\fc;TLg<NJ7&(E6B@#0
0<7Z^5<^e7MN<^ZKO\Y#aEME_2^M,X#YY:IQ#T(6]?^YQHB+.-X88S;1RF-Y/e\?
9J-dKQVd2d#c[aLL47=IX(YTK29ID@1QPR0XLJNK/N3A#LR_7N\D3,AQ,7>)N13^
EU7^gg0&[FdOT[KRJ<)?M56JeY77P0@NbOG,9C&X_E5]^X?&]F09=@9gC73[P=PJ
_>VRH:dF[1F94>XV5MTb)X(CM:.N6(7>=HVRTN\_Sg>S1g,033eG,+:C@4)ZOT+(
WPNA@JRMVI8W-+[+>-9:Tc#[A\9:OFGH6Ug^YH5dO=1Md4c;O^a[g[^?BIDR]3Fb
J8-^J+G/:W8)cMUYGS1L>\W::_<AagV3;L.WZ,]T[8b8E^2C:L&=d[SY>VK;KHW^
,HW0M#NME/c_ALWf^];TL#)0I>CZ2aE:afBYEd-d]?#C,/e\_fLF(]+;[5_SLUU?
+<=E5.]Rc_LT>2@#J9gP?-(P6WO+H1]/Y<=]F<90VHBFUeZcF@SH,>:<]RE]eKT:
1faS\M3UFb(DQOS7QXfSLNgg<8P#EaB^)f#]g7:D?9ROfCX-&R2b.dHMPCa.,<MI
Ub]Y)W7:g.<f,<.P@57H>8JNP(^6Qbg?.de)GeEL6@[_:#\40]QO\I@3?7(^@;7P
A-C#A)21YB5PV,cbJ1P[C.P;M:XAE26fAfeW6@89L=6bbP@e24G;6R_W0@^FBN;6
5:VN9HFa75TgB\faK\#=)-gHO3LLcX&:,^UP=)99TOWRIN,FLN?P+L:6Q[KfW#V-
OKJZe?MLg1STO.aM\L(@fBEb4)N0F,ONDg5#^gXSNFB^V?,H-eH53.Z->6?+E6C;
MeN\(I/=-XcNEV4&(e4<?SB:-)UX_8C#H1+.@(WU]_T?X30_E.,3^TVCZ+8/(fAU
H/R]MOZJ&L+@EF>AQW@2I>[6M0S#,JAffB]:#UJWLBDc?OII[/\I>6:B7ZE_^BO#
T43KWRY#M^K1BM3(S6Yf6O?Abb05C@Y.603JEQb@4=/EDYZI<+=NC7@+0\-dKI[\
V.0H?5MVeNcYM&Je-;;&[KbQS(MT]dT?#8A)MZ-]9L63+7g8A6^3OD1^ZVZ113/0
7fZ4dT.(GBMKW=/CP>3(VaK43]IBOY+I>D;X\TB(UF;)2_+@\Vbd^4FgI98aC@?c
_#L8A8#PYB?K.a:Ef5CZ.JVA:<A-O/OTRQ@;c,Fe7]:\][J4Kf.9>[GR<g@^KHPc
YeHW,=ZXXLL+6O6_@R>DZO;H?963IYI;2;DUQ-TSF,2]VR:d[YOKT97WFEK,B1&C
GQF+^OdV[7f&?N79b7Jce0bUV=L//e(g5aa]aA2]YSKW><[.\,b055E_,1+)=5^U
G@P4e<FNP]5>\a=_8Ie(3gK/44V7^U0E>T54_b[dM]aTHMSI7>_LD.#RY&Df(Qg7
Of^0A,[UKC3,ALQ?(1B4K()4]c/fBIP[cBe@Je(_Y/(5;2KK,d,Ga4Ed7f9H/RbQ
EXGLEF\89VfK=YYWPEV<Bg?>KaHa#4;VMWgZ.f^:K9\H2YWDD8S47bM(dH[7DT0:
0d)6f<)1Tf]2<S]a@fQY\+?UPBb22O#[EZ9P4U,N:\/+2QAI-H1PgQ?ABK&a0#D]
_G5X6P#/_QKe?\&-Tg2+VC7?Dd>_N8[c\CDOR^+4Kb^FN2BXID_N>P,.a4&\O@Pf
3<ZUQd<bAUA2<BDW/gC](KYFb1X]O&LV:,-d?XRBRedXK;D[I5HH5@R(UMF4<GAL
R@a8eGab5J?W=aU\^bY::W,Q+/6V=[X:ZE,0.:^aa45H-2JY[-5-V+D0QF-@=KNc
<D^&:9,Dg4RP/G&J[4Q9N]4fM;H8.C[AXF6:;20IZI-4CAg9BUbRc6-7g3HS,g1b
2AF6DPd.V&0M1YCKJb(.P1&DMVYbH-6,LI0>e/TZ;F8>/1;4.P1Q,M[)PR/\R#g/
;8[+/Ca#<R,d&dQ)Z#c2F-=NDK-(=Da=c,&F0PIZ2W7)bNC;IHSS7/LDSb:1g)3)
78BE4]eOT#aPgL\V,T3K:HQDT;^N&Vg_=VM359OU.VHe<:gWSJG10K+VU&PC6e2Q
;88>Q_U.DaJ/URIJ=A<:bM&-PEM:IbbW.A+IT[)KLQ-F]4_E8E(aN\07?YU&3=CM
b6GJV]NCY])CaVPK8X<a\[9:F/W)8;:1Z^c.1S?=M&HS;+Z:d7b<SO/aZAFA=AJd
C=;,GN>)LXA9(H7&__@C[GQ#+aHg>6bAHeZae:[f[FS6U&ET\>MDK3,@G)H=Gd0c
^)eXIGPcg74JW&5/QB@f^M&8&0acK[_@38-Ja^EXITFOE,+LUb+4(dKNTc)J?UHJ
+K&7Y7<cWO063N\8[^@-L7]feJ-P:BVS,Y>DG+<ITb^\70+P2N39.Z@VN;[M9SZe
R1&XI=K6A;^Z)bU5#([_a?U5=IDa(:ZVHbf(=bD;X2=OTQLWO=?MaI,#?^D]3JF5
\61QP5PXPgX&c>&bTg-@XNC7<BXV^b;&4NfWWU8J[8SI^.VLLf?_X:@YU[J(>:L5
0?H98_4b\V4g/HJ@I9\:94;:[eQ.[M1[=:SAOW<<cRBG(C56dFF+GYRe&MZM(0Ke
A#ULb:ZMOY+c]A@,O)@TE3d)O=8ZR&8<W1G_ZQYN/XR]+KDFc7H3[HZSUa#0>+R-
SW_Z=PB,3^:,&ggOdCE@9e;Y.\?b9Z]5^1A5YASG(173],8M[dDc9T.YO\7_[DNH
(]N]=HY<QOE/]eT[XJ-W;)0f13Q.L]IVg8/dJV)He1[T?29I8IIEZ2I\X(C0D_M]
AaeC,?Z^H^_?[F4V>_fPDK4JEMXKf_<RGIDW..=+OFW/,_#[&=<A2Q^L\g1e24TS
W6F[g-Q/BaHL\IC-acR,(92MX=<=JJ>@=Eg2QeZ?>]Ue68O^d&=ZNB[13:C&QI(Y
gN84__bg\B^\-Q7Q7UTA8ab4,G74.f^c7?(L0V&g+0T?K&OM?F#dK1O8e54O=JFM
7)cJb2d\(D7=]/aLc;g68c\R\aKET]K<5Kf;/CB4X8(1,(;G7R]H<D=SH@(?TfbH
3U0WWV6#^JXQMX-QKJ^BIA0AQBU?AdE._Z0Ib#R9<3fR9W#I4#;7Of?f2E67BO(C
\3GGagQ5)XXE.M?:f8^^V;L,C5aP>@:ZZ?[LEc8g;BHd-G<BZa27EJQ)KZef@-&L
cW.-9B@e(3V3J4B#01].YV/]e-&3f)),&DO5RI<PE)7cc9&/(EXRd;6T,JNP\2S[
Ig\:(.44AXR/8Cece8K48Z(>(N-[b<BcZ?47J8M[/d&I74LQD6_?/V)6VSfFf9):
YOPg>gV5\4f6IFRGW.#^<WIcW/^cIbH.DSR?Df6b<+-Kd3_C34@@1U3L3PQ.?(0H
R^>N.(e?Q2+(J/>FWOd)KP=Wc,\UM)HG^.^VW\[^8J,9<8bI^GH?+4c\D.O7EFY@
9/@T)9WA1L>d^_XFP,/P3YDB?9:F3I=La5]a\J3c2DTbGB/R#:HeVf;B/Ka-1&HW
SGTA71ZY(d>NV=<SXNa1b66RdN:N>V)&2[HF&2W]fb[F6QUP9[gNfQM?_c8@12GU
e&CT@g&V\Z_/O01Nbb&@;]a&=_QM&Ed+5#,S-QaM(@gHeF3&H(OH92(Z4@MOf:&X
?,JV35cK:f=2(#UR#GaX[b7L9+4C07\6[&P,?1<RCBc-)-cHX+K&V<@;\+=_4V?R
c80+-?)IE;;RFQP[@BN(DN?c\O.UWP-_ZP+,AU25^fafS?TS3NUc(J8Q+H[S9#4H
X>U;<#]NSJW^C_][8I(.WE4T0#C6(.2YL845C98H-<b.=N]XD_BZJ(LP,=>D8E7H
OT0T6.R[XPN?L+gJ)RB@,EQO\E-#0=(+.L#F2I(UP0PfXDY^=M0QG7N2&Lc-c;>I
6AZU=#CP?5,?GFO]2#:5TAY(5YV#VX1OGe=XSN.E34UBU23M>?fg@?R-&MT9?^\0
?D^7dIR/&H1Ffg:dRd1LHFDGc@_dV8)NEO+3XLXaD?YHg:_>UH]J1;@48\[YfKTT
eAfQO[3(8^7,P+TCWSHGQ<([Q\.bM&][4CQ/++OQf(<7@1V2Xb/W[J=(c[JFfDb8
d4(?7FED))#;ZNZ@A)=+.^TKL0d.Oe=^;YN4142VZ=79V-AJLINPa&KAbW\G5g,c
E[C2S5f]I8(+@WBARKKVHIT28V)2D5ffQR(03XYJ<2d]2-H=(08I.cJWKDLU4Ve<
XU:RJ1[26.<geI2_P-Ka)eMR>_JBEWC[R@2R<]7/6I@TB.UM21P(2M2WJ5VAX\Cb
EGM8dQKX2N0/cHe;4gUR,]N^#=6]?;&[--d(fZ2(Z4@&:B1R:UEaeUV8OHV\:d.e
<3\(S\H/;:_3g9#gWWRNH,/6-,b8Dc;P2BUc:?8XWc37XaTg7Z-<2=8D/D28>Q7/
a=YP,9B[)b&@QKB6HO267XV<=C3;&^.F/\@4GNPABN&=N4a6U\Rb;2a]dgW;fMXd
C_D.OHF332LJ/+O[88H2A=2]XB9WAE66,LWZQ,+..b]_UVG?OGfbVCMe.;K/96ND
Y.L<fc1K2NK[FdbOM+S1CbbMV)IBF7<_&>g:O21@-.(0b9<A&R_]/><5#0?0OaO&
@CXTPOW9)OYH@G@X:^aagH)(K&_PfaOQ+\+[aIQA3W.gI-B\:\OE271,#aH\0^d=
XX&U_b4eUDH^-3cZaI)PUXeVJ1W9&WB7&1JA<4@96Ic57>6&\Y5#<P=0f846G-A>
5K5G[25PZ,EbVZ&HW_LVTXbBZBV1HUD3PC)bT)g9\\6cDUKUU]ZfXU;Y,H^Q.\.?
ZVZ0?BAg6TN.=6/9>\EQKJ35R#GS?OD)4:b#4=#BE2^W:4BZR>OQe[cP?3D#S-3&
+]D4>gT]>c<7RF2>RZ9bg@HAJJ3ce#-=0fBV7gX&gSgYTa018T]QTc04)b&87d\\
+1]+(.;9P4aBcU+E,];8EVJgIYP+0@;R)A;1@Z^7ba]d/1G<QPe]>0K^G+VcNB.)
eZGE)U/NCE]_373Z@.dTb#c)/;(LK0aa-=UVNII.EVJR?agWI8ZQ8_=)@G6\@Y1)
eB5;4dNNHGJQbP#e:;4.RN<OU,[I?Rd3H;H0-,B+:CGDb,1SF5-:g&gRNEf-WSL@
6INc;@1?GC7=L?N&M?K/E@:Y7f[F-3:LgZ=>0.?6TX@e/<6F=f:)b&UbJH7dI-dB
Lb)Q9:&@N93JAa5Zb]f2UbfOX@V0L<@7aG<M<Ta<:M@PF/LQUSf5T/Y;U>H^Bg\e
^HfJAWZ[NcOb=aV)Q<:@/SG7[2@;AUG[LQa<TB^Z./K54I=Q6BD8c@]D7,Z3aIRK
./.SWWg_W#0>c.a)C:8X7^K1Ka<c:(H^J=@g#RUA(Q:[dc@&/Z(R#UcK[LHI+ACC
,W\IJAI[EZE?HS/RgT(Q,14VGU?A+?,)8=0M;6DdUR+/M4H1PYWIa^=K?RR#W17K
;]+>1[Wa+g[A7&(E>gX3\,Vb#gW(dD<3)F[A=]fTAcP.]EG/ECf)>2_(5S7_?e&8
,4WS2(DR@>D)MNE;@_<E.)WUQbbbOWeH[.G<KBN-8C\;HS[D?=S3>2T>]J4dI_NK
bUV6Mg7E(_b<L2dAXO&4a0-ObJ98?MNZ93T;@],,6d_c<E8XP+bc@[I)/T24VC(I
Q+OF30&,2D<SKR.g_S2;77@cH_D51ZEE[4[a:?F_,#geFY3Wf)6]M9W?IH[ZQ^1A
XgHgbEF\O[L.]5d<\=:3^(KK:Z^RHe.[D2a@6,/&[P?)&KNJLe=YbI_EG=D9c&^F
?JM52?fZB@P5]bMHgIEc,@JOd0(AD?c94.>2/(bK;[Q?^\]>#9R9RU)GMfHVgIfD
5I:<@E#N?D)C>@R[S-gbH@WFcH,aXc\d:NN^;Ge7VM7D/K^[T^M#8YJZe/)N?\CZ
S+,BZD,PP[6=G_87OZ2AKO[623OIZ#<+X0/6^)1Rd_TC&)0Efe-<M/FI6eaFNTfP
/ST_bQP7S1_KaU#TRR1[^GZZRXJ/B3J=\5>^9>XHIFB8B/)ACNYMAL9,NLTUaUJ-
R>=;D2Q&5/J1G8H<IO\KNHM9-M==C/_<A2(A02_RF>VM@eUA)dSd7TYg@IB4>88f
AVd9OW,B8,1BdCOeO](/VABTbFa2C^PWfO6c02-Qa]5R&+?\\f[O3;M<AILI)#_Q
JdL.9ae^bgWYJ-7g_2846Y4E3=3\+08P>K[2BV&LKe+=(ea<I\0cN7-+\K9e\d0M
3HVR4cAcHDQBa;6@U-ba],\?E5R@R1P+]68DD)35f0g<B^fLIVEZdE4CL7^>R+QD
9)V6U<.U6=H\X9Va^Y_TFT0dSac)1O)(CYNVb4XHMb\(OeE_L=85\>cL)G)LTD]N
8[JHISAA:BY5WE>0f@CR_(:HO9?#DK]KY/?E,J?.FAc3]eg1FeN62851d-])HN3e
)DcGD)/7MGd;&,2<@?IB/Na_ZKGH7Cb8?2J+C8Fcd;AaTfa3eR)b>D5EDG7gVg;4
V4)MGa_3+AOaL<Fb77_:0^ZZH?aV?[ACNTCOCMg8+;02g711DHScZ8G<KEFgPOX8
)1WX_UO[A,.#-=[MSYb#N=g6(LV8Of(NA_3),DC:P0UR38?OPbD13F.Pgg3W?9V7
QHY&c?>9V:>D#&]Y1c4fU\]X:8.33=)HX<(V/9gXMBe=A)f(I)U&bW3BX.e;.3FV
27/-:=>L#5VD^+,/CJ+[,UO@[_MJ#e>\QA0A6WR.9&7+P[(8K]?F\/H4gAGK5[9+
[K7,6DXgG+(9gM3SXR=_^Bb_fJ-4<=ZQ:U07WS6?gQLE(<A49]Y5:gb>LB7TP2PE
:9;?VZK2_W6:CH&,B_SCXZT?YFNb=7J1QXcI8JaFd<Z6>,\c-QN9Y:2WR(JOMS.N
Kc(]He9,--\TX5(gJ:VE5)3?;P;2?(>W@BLNS,e5C]1NPU[cRW(TS2H=,<\c-OG[
@cGS#&ZeIF\X.BJ@IHTBXBW37KTXVZQN35K&=^8KJP.c/:ALT^/D4[bG\5bc-0#V
:Y4CS3aJPaG#I[>&9A^ebdUU_6C])bJA9H;[edT^I,dQ_:eVEF#T@B\/g+d\Ua3G
GS.EW>a?fZ)F_Kb1CM7Z5e(2BC<6dYJa2RA;QS6E1UA7/03Y[dXTY1^^Fg?YgM<^
O/PG)Q3da^BS0J:9\a7d#6&8>\(>E<#\.H)@,7LL/RO]bMC;1FFb1;aE(0XZ([=A
2Dg4_0a<53AaCM<)/L_gQcV.VK;a;49#dMNILdEK;HbgLJUXRWecbTVTO9ORb_eU
=HKS1faXL4<COaU^MJ_7PJb:g[c(9=4.+caA+.Le4&+^4Wd<Z\c:<<Qc/R_Y/@NF
3dIY6,B7+7+J)1\5K5I.DbC,a=^bXJRa#4,>^E7@>dcZg>LeFb=?<RNW)\f0H5;]
IN/HQdID(gYBJ<S<bNLbaD2#WV:Jd84C6@ILPLG,23=eWWXA:c=I?K9K/\XJ]YQP
?)eVIeRD7&2d>0A.#:Ue&.<aP)e4-@Ld[G6DVU(4b.C,MO(g>D;a53V]9>;Xe<1(
L<22BL;?C3L=/b]YQH/OCaRRW\7Q4SE;VSNP]609.41V.QWZ#)>ST?YGd+SXG(BV
0+1-&A9IbaE]AaUe;OQ<AA@9OA_ZOd;Q[?K5Z-(#)NC_O?R+H+=fK</DN+WT[/O^
P\5@NSONdWaCFJ8@Q>@QGL#80A.,OP<>]KKN-J[Gc\>+ZCT>&N4BNS04:=^/Q@a:
bOdVLW,Q>(7807;)S@H1QG1f=CT<0>1?+(B&F[]0dc3aWE;KR(JU:<.g:/IA(.3/
C)//RcaERHQ\=>([MXAaTG)BXEW+V@9<LPSINQT#;TZ4]^fd3-O0fIDHT/>QXEE)
CL?MZA-Qb(B;G/gFF0.T:#R_dB>]FZQC4OQW7N;DXQe0=/+SK;(gH+_D=@:.GY\\
UL3/F?a/M]C7&Fc47;[X5ce7ZeR9[]e#>/A]Ta0;^MLTOgKTIVMVMBc<e[UF[&EN
FH<^GOgBEMY8Gf7P^8MOM?ICX)NX#F6(.S+B(NdK9a_XTP^afWgdT1JRN:-f7K?S
P(-R]:dATALVCdWd@SCE85B23;)>TE)<S#0DNM7/#Z]UaZV4:B/F:RA6-89,@[-T
?JBM,MPZ4(Y5RF>f5(HV#9BS<.(Ja#AZb@Iee[(9S6<>g]a,Mea.gY<0MC(9UB;)
WbOO&95:(H&(b+bRgGP3RgbL^/JdCDX6_TT,-TdeaGF9XECc6OZ^?+T23/CBJCLJ
4IYC;A4Na3:JF#?DU)9EK7+R\-<H?[-W-^TU@&.2@WSa]b9fU=1I.DVO(e5.?T]V
ZCgb<\RYE0=/89aY5UV4#,P53f#\2FV8\GALf(ST-\J?SJbG+LR/PYPQEFJ@dd8g
ZHK&CO4\,MGG.1L3I:[(3XDQ:DR@03RB4)^(4\IJe<bVXDNJJ(Y2(aL^I=A(KMZ4
UQ5-0<_=M3/39_(8T<fSM9^=;?8-9Na2e_2GKaee9PI+^Ca7bUf(;/9#Bg8FYW7L
744.dE-MdXA3)4g7bOKFPRB4ND[XeU/Z+OL#[Z+]A<L[3.<bI0>DANcGMYV?6./T
[9Q(Dc3Fd;+7TAM+63H\g>8=)3Q7b0EO6S6.6@KK2dW)0.FacMg-4:\c@Xa:TVXN
FICeU6PS)BU_A,>ZIOS3@WWQ[3b&&@O8W.GbX+V=X5(#SU\I54D:(PeOe[J68e3O
\F/QgK2ZR&Ud@f^E12.;ZQS6SUb7d.3B:X,-#II@?VMZ/J6?[37=;TNOY[L(0U2E
M?&BHf8^W(dCM^&^QBW\Xg._054D,:UCQ@ZP:B@F.3T_bH[IOG.V+(>F1<Be-6).
\IcV\=5.?LOM4EV&?E?bNVXcLU)_c^3+c4(:-(2LM>U^H2W:d#A?E->+1ALa0;4=
\UXU]L]0cQE&^LLT6W=OP)O9F[<KUE5d4(]#U6_C=&^(?F)aKc=[&PNK4Bf.&(M7
?3T:VD-RM><HCT3ZTAD;<UfCYdG05@.B2d65H4K)LCX?>McNV34K\JD-VDGV?A4a
<P<U4^VN&Tc;JKaKU:X#YG,:c1;O1HS\7g0Fdg,S]TJb^->L8>8MK3RZ]2fA2KG5
N(FbMN5^;#6+<LV4BZ@2&>:EU@;R\)fDMUX23^];AJS+d^ZQ@)[;2J1D.B,SE7AF
ggdMS0P,Z^UM6g/67M1X,=8(dM+>(UDK_\UM+<V(5@B/>D;RP-Ad1QM/4]P&,]6C
c+32CU^H<(T,@Tc7T)(:?-MV9I3#H7V]C9SI52F9E&fR#6CLQ&KJL=aaQ-&9JVd1
T,#&W6:X9W;?]/U7<GJS^cc/0[VLU,C>9X=,VA;<Cdd]b\?e)\=AB=Nb6G&.CX-_
SV>dBd#6B]5YR=7<?eN,0O&6L3Q_KUD2b.d.VDcN9]AFAEf+4FD[#LSY_,gX2WT-
./0+EW&d>)5b+f7U_WZ:Zc#=Wdg_EHR)@\@a)?ba]UB),=\3dRg5I.=QAg0>AL+?
FUc,9IIK10Z>47]e^_P/.6KDCXN#\HG0J5PFgHDHBBd1YTXY\0]/#cB/&B=OI6Cf
\GYANYU7a:WP3#D6Rg[O1RL]\c2>Z<N9[AMFT5KI44I;9Ae;Y:.BJ0bMLF5Z8CAV
a1=CH9>f:c7=:fAf-<;4T:g7<:W?>Y4R9a:YN^PbZUa,,X.\gO0cGC,,-YH+M[IX
bN-b[93Y?]N^BV3H5_:S)8Ia];c;0XEV](.6.82>H_bB,-1+5;5P,#:K8d93[H4B
_@.A9b]GE0(JbPeaWQ>#@YJMHDG]3DML8ZCJ;<FPMQ2-]UM(0M]IJ<E-WY]=4g-A
V3\b0D.32cKMR8P0FI<958P3AE5FCdKBB,<?b@e\VIPccOCRKCJ+NbN95MI(WNQg
ed^/g,GR5O=[@78d[Z(@#.J(L,0^_PX>8Pa;,80)09+B.T^=@)?V@THd6a8#]Lc-
4MMM4LM:^\WF835U<I.R8P+=,f=>9S;eMET/eF&AVT#C<B^8)cbWUdc)fCeO_DM=
NU7R6##-#WJ=#W@>7<&XADeC519-)4J&&a#5Fd?#QNB.\I8H+.?7T]EgIE&0<3=)
\^=1SX5g)^&?T.,f4?IgWD9QR_.c==L#cG=.;9(J0aOc#>:VBT/,Td1[(EHT_YL@
GER;R?N]),,S23UFMbg_2PQ5^c6bb+f8(6dZZHa+GZ^08#Z)KH6g3TJ853)QE(M2
7=4GPR@]a<BEKN@U.>FJI;f>##E./-]<3H<,6VbB@?bE/TW6M=BJ]U#J<M&IV=R/
efV&[-9<S_d)&UZNYD,9GCG;8V7BT>)>T]3(&Nd338).S[e_-I2SL#6DR&/ZD:H?
40bXegQYNV:;J)PY-<XaQg\>=_(H?GQ+;8370Y+8AgI(U(]WBFPZe<X&./(=F5@W
M\>Ec@WFKdIX4Ff3g&fA@Y?KcJO=L\/EGFU9O5F20HYUF2)06b1^#&0K_2,HNPGT
HZZ]OD<JWNI\U1U);aW.8U6ggfR8_cf,D1D:YP=:SYHD@]RdZS-7\&ZL>_T_C/7K
Sa8QHMTD[6da#BI_+PF9.+VHfG&YcJ2(fN9Y@6ZHfVXZZNX.V3Vff8IPV_L\UCUf
5E_G[P\>Id3&\(A;K=D3>2TbfW[eJ#.:MXLZ?QIb-GZUOa1Ug(26dHDU6X:\)R)5
CM?BV+X)Z&K0/3^d27>F(Y<U?SWCW)7]5+a,BI&R[8d^Me]_BHAUY6PWDMM=CGG>
VgNZ>^MI1b:<?Ue&6FXf+daE==&,>7^+7FWPPV^#XG/:)1,1LE9<Y\)E?b.YAXL^
cY764QMg5T6cZdSb(,/e309Z9?[7+[FDBc;I6#=14^LQ7ZLRfOZ(X+[R@Y-;L>&I
F<DC703YZQ0/I5O&XA7C>?P:6f4&X;IX5-(e=GdZaBC-9Tc3DL=C:?7b;-bJPYeL
cYN;P&0XIaggEb-X#T5/[H[UE10^UM9)6Y[c2@6fD==2/H&P,^-CHE=eQ59U2Z<e
NF9JVMXSEJIO4@1T5aE/>C<[C[Fb7e=I5:CU2dB-]9&;RY[;E,W:NB(cOUP&X4dA
\XO&\ecG-2@.M3<023FZ^3X.1)7EX\\BDFT_KY_6(gH[56.]X1#5/B\7S+1QFFG@
:gF<05D>#BgR&).:SZdRVeM;-7RU>C5KN&S;g(YDO2W?[Y4c(OW-X9SPH(QI<-\b
+3>f0O,De)fKF09a;]V1TC(GYeCOCFPg.UKO+6fQ=8UQO-27)@2I@2g=K<RbfU-;
&VHY,]QC]Ab0XL395#2M&CNO=L0<?cS3P#::KRb.H]K=#I5Z._W:,=,O<\2A&8bb
8MOR&Z_T;e)gJR_NKHK(;#W#<PL/HH8d>V?P-M<?]<dY96:8KDH8:2WTb=c##\=D
&E=0CL9KBC0^_T@_&TO&:AGV2bO0K/FF9^3JS:M/N9^G;(;Z,\4QU):ad_(Q?GRG
#1]c5;=2;4TG>aHU5P?S-81XOIOfVPY+_d,XRUd<XF+IQ#+C3+)TWd86)\.#IC;W
a\ZQVcIZKfc:;ET,8gU#Y<+6Y+U)ZGe[&S2C[33-+Tc9M:MK9)g\VN59#R@[&IbG
fF_ce+YAL;QRfcdRfN8d-1J@DLF7EU0g@a@WfOOA(P@8c9(Y]J4)RegY1Lb4C<;C
((Q3W(8>@?>MZNGAe9VZP@Y<d9GX)d.[ec/]V0RP;L5:-<HBePPN4gVX\6T1J;:)
;Z]1f97G4H>@ZX\^d:LD.gHQ^XF61Ld>\3UbYdP2&DG\#F?ff\4WG2W_U+g1KL4(
\?_DRO+,X>4M91Qaa9^cdAP^EAe7=O6H:;/Q)R;GaA63N\eZbA;g2ILR7E#NI-c4
aF1aaR]LU?NMUYQ@96ZAJgYVM@R+Y9=O],UM\f65;??(\?\>6L-5-E#P#9?M(-K/
4ffCCYKHO-aKEcJ9b;FUfZOF>G3)<FP_:L3;=Q,K),=NeF,Ne3Y,NdCS=OUa=:W1
BQb5O3MJ<BOT9f<=DK:dU1N5^(8K1OC[.d+.U/Z9>gQD8A6PNW?dA(/H.B.04W-c
8_:X+5HV9.#RZEB=&dYWA#3<gSUXMO]RHHAYB;FCGII(ULbJ3c-^a\[5&_Ig_ZX1
>.>E(^\b)[M(?X7RMODX#;gfTAN&PFL#O<.eAH^OYU#)d@4DAP81,K21WD6eIEV#
752<^(Z/NfGXV&PY-B068dVD@#-L^8Z6Ig9Z]2UBMZKH(]OY1deU\W#[4BZR^O[M
Z21+gIOX@UIVUV89M4;6+(bE1bWfY[\A+@\H<PT1.64A#DZc_P.?7I>=?T9(;Nad
Za-#aO^8+I4>B21BPDSc6BFRP,H2Eed):$
`endprotected
endmodule
