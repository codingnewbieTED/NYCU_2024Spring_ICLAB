//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2024 ICLAB Spring Course
//   Lab11      : SNN
//   Author     : ZONG-RUI CAO
//   File       : PATTERN.v (w/ CG, cg_en = 1)
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   DESCRIPTION: 2024 Spring IC Lab / Exercise Lab11 / SNN
//   Release version : v1.0 (Release Date: May-2024)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`define CYCLE_TIME   15
`define MAX_CYCLE  1000
`define SEED       2024
`define CG_EN         1
`define DEBUG         0

`ifdef RTL
	`define PAT_NUM    	5000
`elsif GATE
	`define PAT_NUM    	100
`endif

module PATTERN
`protected
T]F^O0F.:;7c&I)=@^UK,Xb@.MRe46Bca0[/V^M.c,6O1MK6GQ8R3)/&U\dXa>TQ
]c-ERTYTa:Z?ECIK;ag)#DgSL/]b7.D9Kb)EeV[G0Y1.13<\06QQ+BbL<bV<NXeX
d2\7I+?A&+GV>-OBFf=\GZ6+)+P>,4]D-[L#O:R-c+XN>C3OZDdScJa7PORB9#KU
RR,14&6&K0X^d^2MPPRY0GJ-[W-#^3gZ<-^:D8T9EGR<?Y52SdS<0Q]2aAVV3>\d
c+PYIdX>Lb70B0P0F0#M3;T^S5?e/0P0cd[(MB\g#OMJ[)5R9VXJ>;a8EAgL@aag
;^)@<E.eTPD5;=ES#&(f&PZOdIa+L;;TT^S5[3O;,NV>_=PW[d)_@+,2A_0YI#1#
;B\]L<GO;+fRC=930A^[E)F49a]0)W1dHeFYQ7N&a6e:b+)_a8W@a[@gXD.e_JRQ
AG3PH,\f,B,D4.^?]?KC717/V[g_)(BM12@#6f0@XXW,c[e^VK7#-7,0&c]7=XNH
Y5?I0J8J]>(73Y\15+SdU,U3cTXgWIPHQENS\;?S93)WJLD_7[Jc@U_^VEOIL1DS
YM\^[Z;RE^<UUE;L10ZQ,=T=/W;NNdC6C:);23B3A)gd5aU-L<+-\RZL-I[>56PK
_-4F=2A=Y<J3CR(cWB:NJQ7?D#:P(DZ#5d@Ha)ESWFI[7S32RA&TD/>T-ZWXg5WL
4^9C6]?\_NV3X--]1P]T;H:JH6UGE^5R>G^e3OB)#A7B#T[A@(a\MG,Qg23>LV:(
V=@cf>U)=2>.Q#+J&)YA)_2KUJ;E:[Vf5@cT?1YD3(D_4E/W\;gXVI,P95.HR3a)
eYO@_L82cZ6e[&,=6-Y[gW&g=VAOU6;.gB3@LZ-V5D+Gf3E>.LX@,BecS.Q(a.-]
/RafX3Db&Q]Oa:/Tc]N^[b1?5:#.T0?&#agFX79/N#W+;H=WP)8@-EaX?]1#:A[A
2LGLK0GZB(+;<>UT;))aVd(4G[7>TG?819,@O]cNAb+\K_B5]8&4ATCZ@]5V,\\T
0\Ie(OUaSLY7eC>dV:ABb92BU\UX=&e)6Xc/K+GL:I+686H9OU4B@gS[BOVc8,9<
6X_P3OVH4,8FDS5ZNdMbNbN22UXZ_7?WgDAg]\;HNb4#&ESV1EMdO#3R\6]BS#\]
beRW^fT?MY0DGO:JVa9R^J@Fb@BE,5WaY\++b?#((Q=0>Rd[>aBH1WSWG<eF_FX5
8WX_/7gACg\>ILg+:+,;T6?BeD0gXIa:QdL<K]Oe4_NIgYf\;-Z>L&e(F9.FbB3;
JTU^fg05SXX-A/T-;@QQQbJTD2<2aa83Qd6cBgVYC4..4d^YR#^g8A:#Dg&YBd\8
O,U>2[2/GaJS0OLc2.CFHQ5Q6W/\KdJg-QdHVK=S-ff<c+feOW;S]4)O1gGY?&OS
XA]SaaMH5RbIU\EIO?6K536R_fTC/VK./>f(TR^?753?=V#UN4Kb3)R7;Q6;\R_H
CF)Nf_d?b+IXb]?2fGgUP]G8,O/1F5LNLCBUa7cgWKGVLZO1_X?PN/KVe7>+fY.T
=3+;A_HB>-[c_=K#;<CVXO[9+1NT(5>R&Bc.\SJ0a18US5B.@P#(),cUdbPXWef6
&#=1&2O=Q8@8;?RWOC&N7T1HZ+WXZ93@gI/8<C:cbXPR;4)a&)#5W@4?_^WE(?V>
e6J>1edK_ce3Z6f9[&,dE1JOX5bBe]:NVWDWY@3-HY9V/E8QMGP85:T)-FKXHJLE
B32&J1G+B/KPbS.-7>N7.6@>4-5b/1)VOc)J<[^b=F64>IS6Je65A:8K[][@(QRF
^[XB#gPJ1CTA/8FVg;?g0CV.0]W:cM\Q;U[?A/#AfDP+)UVHN=Y)ZSK_c#7(:V?/
@E46<fGMWVVFSfQPA6V=CFb68PDf-PI@f+8E0SUO6CSI+7(FGFJ18.W<>fWD&[=U
>ga6IR2V0>#&\Y2KZ3c1^];A-\[CgKL]7A/bYY@/FPI.TQK?3f5PYK9-C&1H#FeY
HLeUW/b1N&V25fM\O6?F#D80g;W<Wdb5HP_d[8[7+Y&AXa>,bP\)-^M)FV:]&bD#
^gC._J78ZM@6)06<YYBO@09:Tf2EdICFa+-RT;OO5+O8S3),7_J[I[Cgdc\]FF)L
Rd#e(:FETR;^ddU7#W&a&.YA-U)G:^:L+20I@BT9507=+/E:gBGUf3W/0J@OgPY&
ITA&C5KLG<e8e,(S<_a5BT;3LKfVcD=SS08<c)PNPcMUX4&_9_7)4-Y,6H_/IZ9?
@_&ECF0f^3MJf)<d=UPP+aSD4[\G>N)SS5Wg&P&4e;HD&W/1@W)fQ?>>a<RSJgTS
\,RMP>GgaJ,@#I7LV#1EG_c)J)QBbA)#_0dIRa-4A1HI?E3U=K7eTg4I4a&b@9[>
27L>I)6cU+6.<^COgW3[JL?Q2&#-/67>](^)L+H@S5@@9H8:22V\C1]=fH<EGa=S
45E[d37I&]If7D0ZT.5/2;2]O3CC81<6,/2cTG=]U,I.4+7JR1;Xf2bR#V1=D:OU
,Pd^SI[QOIb?@Feg.U-;EC.FP<BQ\&a>CGY;dBIVBLO1U/A,/FUNW@/86N/Y^a^R
gA-[)4Qa82:KK\O+f@+(U#?YS5#FgMV<L<K1?4S:/U6@TL2[S_>Q,/U+ggPAD><R
;befbe+(AMXKVdF6W:](C>Wg9f2./[QeBWcWSQ3())bT49ROTEC+(5cQH/Y5N220
NAf&c3gE-&.&J:,#1U&R]M5I&LTWBMD+,cGdFK>.]Y8,D&WDD32&f+AdF+_S07\A
9;Q3^=V7+&a<bdJ66:NT,Cd1<(RVg/gONaZ8_6_KIYI>ZR=c@I=PTOWDDAUbZ\SL
;gPP6;JCARX03N>2T<#.YVSc]4c=cY#V2O#CcD_ZTab7[fWRfVZC5U9^g#@/@Y=[
b&F7-1=/IF8;<4KgPQZKC1<^1^;0Y(dc6&aa27Z3b.6AL^4KOc+7[1c-#f#;\BOY
NR[Z5+OSY/6R-C;:)A>,]<?[6FQ,[)ARW41[&cGTVH)7DA>/N;26XVT2[fY)[eYU
T(P-G;/KLHT2]:DTFcAW#TJEQDe^2:1(BWggOPFN9L[DedA48b09@VM3_2UdF=+K
_Z/da+5eT=I]YSa@5[-\]6I+O7=?MMaL.N1E[2>;DYDQc]2KSWgDO<)5+JQ#2350
@8W#Y5FT-;;d2P/&U1<0N82N&Dc8:[B2JTL,A=C8-&+,Z9Jcg\6Q2;J66RB[ReU_
/fJH_BIJD3Ug#Y4SVMaN,2.Y1@9V_XB145a?L-=<ONSX5QYDcJ=OQ;3MAGeV6gZf
O@;KBCB1SWFV6B#E&a)-OUa9^aEP?GAV^d/X_(LbJJVfDd&@&^gQX\PS/AcCZ\SW
31cc9&d(EF\9#C>T:#1<>F[&YdVMOROP>FBEA+2fMIR3DL0^6YD2:=]LD)3C/P)&
F5?5SMEXe7.d1R0eSVA8_3Re<eI2XYa#-dIUP]=Z(M39R1[F4;)5?UTcBT#C74VI
.AUG7AIWFWH#6Mc\?EVLXb&4/aeQGFeKd>aCU:\g(#1;cb,g;Y1^O^I;F=RF[2[Z
;?g^GLGQeK?fUOW\=+;]J>2I-O/]c3(X35RO-H@O&Nb52ST>+)\;2>6X&gB-?\/:
[S[2=H+VLQRBY80QVPP)A0@]QOI(cb<23&Y?9H3)SEF[gUV[b0=+G@eWX5T]-/Y&
/_ADNfYYQ;&,_KP/0F-JDN@V^)faJc66AU3e:Ydad84OSFFb7Y9g]3be,ZFGWUWE
(JE067VVA^?)]WF392&8+.JO<0ICBb15Pfd.C^&(?92Fb-4QF_1ALX/.:R68dERA
-R[S<-6AR<Nd^b)=U[8f)GbP3d2@]THZ[Ke<Z=5Gcae<J:/[=80]a66Rfe8PAA5g
^J=S1B3OGKcRQL/R(0DBR@QCUbV,U_129WMaKKeAK;eaNA8&L0L<\MP?2B?:6<eb
e0K2<):MEcU/D/TcFR+O@8TL)b\X.dP9S\X=K(3KWb9BI?d6\,NP6;Y;K).DFfX(
)cgF#@W9[Q:2Z0\aXT]G+T+b5)E^#ZZaN,:HYd-QJ^bWG4@A1d(D9<G#b;Sf^/KC
e&J@73]R[)E_G<>I>_5&VFARd5;M3Kg,)V1-G;E^:ZNF6^T.-APD4)4Y#Z_ZHVK(
H@+fXKO#:5U2NWBKgcE/c6N2P&RW>1W9BNTL[0ObeIR[PQ-R\)cW6g[c\D\[U510
@0,JVP4TFU_#U50cM?G36Z1.&O./27H2QSPB)P9C4=NaaC:4NS?KWS61;4^MRHRd
,MIOe.=VX\daS<O5^[bg=aTa)(?@DG3gb1G[9XB8a@\J@PTO]E:X140c,Z7f81[d
&#d/VYaHCGgZ?;e,[D8LGUBLQ]/WZ)FUVT=8L3T#b1A88IZb;bL8SJ518M&->_JW
MUdf]LTde-cXBFcL25aOegNcB1P=a@L\-T7K2N=>)NGIL+9K<+_GMP6NIYZ&1e><
(d_d]-BBBB0g-ba@R/L,&],[]M(7-.J@SJ4\BbY+5/OZ)HV##.YSeadGGHg&JbQ,
&3?f/>2gA:0E;316W+RHK#27(QDB5[L^QGS.@#&-/LH,RDMX+)]@1.=BS9d_<gZb
K0(>+^+EeX^fK,HJZ7L>Z;#6=XHNB14.,/:GP5-(RKALA>]^AM^#a/9@f-F9:+;&
[ML,[4J7d@9JT..O>&096:)VF,,4<D1GMTZM:dg3T>V:QTI4OV8\FQ9NcDP?_=da
?<D;9]6DM0bMQ]fOR8NX,NE4Q?N/?BA@b=g/U-5:L)<1KOg7T#([02=AH[;]=B=#
SMFa[8WaHcW+[@F^_[NK\(@<RKE99WHMWD.C\;(aK<T;b6G<=?YU)b8Bf:UBY\X=
;L^a\Ee#&YGb7fL[Z91.#?;6XQSM;-:WLEHEOJ1<c<P@Pd5=&_ODaKQ2+\^HJEdB
<R5;W+1/14>1-/?.PNB9.02B&OUQ:c6D@c;2\XS/5;,g:EgH2H/F6(/&M0+QWX@#
)2-M^g/#^S(\,JQ<E)O@:O>)_QUbCBfUC=LF;<J<,C3=N9NUfaLEO&,)7[bU?4O(
Db3AP33@:JVGLc1f<GI3eL2UP:]#R<.#.Eb^217(R)]OT.ING#2_QA8G8_IbYdIP
#G6]&,RL)<[81Ce5M+EAg4dTbJ<Q==L<bS9J\1d36(.fN75>H=W_J434V=Ka>[-&
A5.(]XJ;L=HFN:-6]VR6Z;Y720]UBIFC;FUCW>QMb9J8c+NA4=R-4?-C0bJ)RA,I
NVecQBDNLA95I46](<3F#(Q@A,HNHIQc3J;KGRe,+LP.D9F)#\5DJN3cD<BZP.TI
3gWTOF,\N4E9:3OB/7EbE([gGIM#Eg^X9TP2d/()CW/1Ta,4\0;A3-L,V^(,_;fe
8[d(VZT=.0F5JD];-H>:DTd=&.8a?]2fAIA:Z>G)Z[?M5;WcDSQ408VE2_TCYZ[3
^b>e@(.IJ=S5&X6e:,??N)GO16X2U<YE#g.^&>?bM\LO:&(W.+F?40g<@[0@61X4
W<CE6L_S;^E?g9=&#]&7b6.>WDI>1FHcQV9ZYI23TEcP9f_TDXXY(\L>/:I>47Y)
P\WE>fYa?,RP>N04+(Z=X1>T>#(fA8--A+5_LB=[a(/20A_L8c04()Kb8>Lg4;\-
ES6e=<@U<<I9V37:@&eS&_Q8R4W5gEGZ<c2aJ,d:0(\NMK.S9D3@R[g4-RdW8fbV
dA3;OOK09eYg<DJXY3I&.?K^EF[KZPKA>Z3\A<?Yg,>/(32O#^gfU]>-?XD#P=PJ
B4Y8N]OREBT\^FP.44UVM^[F)GQ3XTZKYD@AE,\)Y]R?LEEG8VbEKce_b,U<B/?6
(K0_Ifdd_^O1=:P]W>.9#[D8,38Ofc5,\)1#18]VVd)3QL+^,T+C\a2UQX,dP+a.
<RM9Z[M.KD8OQ9[YbWW(3W:Y^=^4T^:RbV,;)T,E1I\[Jf)5dNOA@C5[Y;fBd,f5
^9E4:dgVe[T]>TOdZK=c)U)^?<&F0Z?C.(<#R)bP0>^(Gd5CdDeC4;/ae>\70cdO
]4(-?/:S:@Q])d#Y:32=DN:+_?,feZReALW^CUaE<1<DbacREg&aA4(QGRYSG1QY
eBDP)f/b)\W,I>SZc:(d@7=XObF.dJVE=6ag:TMfSa=9M9Q.E]F\+=W:N88=IgD[
O;#,+Z_E5E[=#bT<_QP)CJV2JI0)P3:HSDSg+eLHXU3Md0:gcCGf#&_Z2eBBd-_J
/fRcU-1B)(5Q/2b(X&]eK5APf1gLOGNdg3e&(M)VQ1=C^</T7YB;HcVF\cXMN]?a
4AP<Y+VeD]__4,G>eD+N,DI4/3FfYI(.25.ac3/M+^0^Qe9DMEKc/33JIgW?J@TF
gVF@(MU:QS\2aOYPNJW93C]KU4QF6<#^a6KGL=AT08<.6MM]B;TX#IQE0EeN&#7X
+A\Wa-H4G]7HF)X/\5]E?[e<:AX;D9:(?R.IbRGK,FO3:VgB(Bf>eNg9A1eI96-B
JVASZg8T0Y@.292\ee-Q+F8cf^9X\HV:c6^LE^39FHO+)81B2Md^DKB1-/S2&ZOU
Q7LcX^Le\(Z:4E[1Ra6,+NeSQ]6b/=6Wa>&ZJCFe--K&Tga4W:(INdf[:-Z)_A73
O7FV;I7,.c)<<XDZ/JI^cVS2VC#:E^8^@2B.WO\=&0I49=fBVfZ2W;469>4_VF]\
[KQ-<f=^@.&BXUQ9DYKd0WEK_B/a.0V?FKWESHD&Z_3:U=EdC0Lg-.B.a(cYbZ/5
J2FYKE^6YQ9-&eRB,gO_YV.Z(A6\2Bb[]/E:.PbB>^)+F,MX/&CG?C6;Z\,0OgB#
d)X&f24B&W9(.^H<;a3[^Dg4]PQTP7Pa..aRA?7PYT&d2_HL[2=e<>0L&^81fNBQ
Y69B-(+?fYCQ<LU?2cVG:VH:Y5NBg@UAad>^UM6<X&W/cL_GTbQFO&K=@eT1_&3L
RGG&L+I<N@f07IUKCGg@1<-8LG)D1WK_.:2G8dc_L_5+GF,b1V<fIM6&PSPT8EJ)
(GLe9@?g#KDOZWE)ZQ0./\X#]D&]=[72297@LBB@,I(UOagSVTdY_ac:]5A<#XfJ
@^):P]BX:,GLg2Ec]abYW[N)2><H>b0V):\H27eV3I6?JOS#faS>+DXKUQ\MB0?&
7@Ed;@IgAPfULIcbf2RZ5cX&Se+\+-G)R3Z5,Y]#CTgbfZQ8K7HNJRG15NcFV+M#
74HNY6U0ff#-6/8]>?;L\IeR+]\AFZb:4R@J7\dP\Q/,0,5GHL#Q.;KT2VI3=\R7
9@JZOZ&AOOH[B2^P9F+LK+<VI[-^;,/^),O:+K[CDX5V[7WD>b1gP:XVV=PUgIIJ
^]ZP7:-1,0:CPD9ONWaD?DNRY7JP38^a(=)2<86KeK36dHC?6-+UWEB[O]Z//eS3
I)^K?IY<MXNA0=JQ,F_^)QA4-_D8^M)GW-gZ6/=Rc,;-F4<IE<H2GM+/fMLcc8\\
[CA]TUD5[_M>GK_SgP\,3AaX.IV8<@3N8-@^2dZ48KG#2Q\P&JIBQ#&)a-0[F]bP
DVXRd((B2\_LV\9O=CV=)+BS]OTSLI;VYPc/HJ=67YP-_gg=Ed94K-/2^XUdL6fC
(N12^NXL7A@aAKW&]UX\\BYA9L>_;S].E0P58KC,#KLJ]V_Y2=9Y(6Sg)BRc/RW6
J7ae<<]]2[GQL)8>=NYNeB0V)[-AR]:K0.Ff2[Y.^>GIWR9/Gd5\>@C80d.THB:-
C5g6::6@ege;E\ZT&a/C_PXVdWDH1U],E#?&-Odc)=542E+26M\?PSe.A]UJ8X3,
<=SL_GPP(bc(WK+0V\KZJ74]RKM^SU_Mg1/T.eP;)(?(<C+;g0R-UD?@YJ.[3?CS
HeR;,39fK7AE+9BF^5:H[E1\;f]7e],4[>Y?/[EMSE^,_/AL<RTd\[eYf.cX2C)M
=A#B(XBOc+<PI^O<FeeX)W^7_GVN)NF989e\<d]Ig8KUJ&DO&X4[8<.SUSdX#Z_e
f6.LL8@,&@M/46YW)3aV[GG+GLM<Y,TaQ-.CMPE((XJC&E_^E]@Z/QC#eAB@aaAX
#69US[Ba?##.Z5Q[<UY8-=HO::5ac0HWcc1dF;dS\)K3(78I]?JV->+[W8061L?X
5T,#B^<gD+^J7@0;]Hd)HK78V&@a(5d)W87GTOXgGPcV\2HI2=V>#,e-EFM&\3_)
17PG=f#XGAL5/)dSU]-_JK>bcGbJ3&W^ONIC+ZQJ7<WEVDOeFe&-+[gC8BHJ(PaC
3<(N^(F5-:Q2M&?BLY_T(7d;PUSW#T7-,Q.OI^fXOS-QOH-<CKIDf/_UXFaRZSQ\
>8eLEK[B<HC7,5YUV;IS;JWVaT])U:1N=[MG^PFG]YVCA/#f&T8VNfe]PABR25)A
GPT.BfPB6Q@3VB[H)e5bVK4K51&]+HD#d9adW1;@e/Tg0H;//C5RE7H.9(@U81E#
V+,,[Ze3]GBU,_N./9S_&#;fe?cfY;e/C(bebLAIK0SVfM,>,)cPRMMVa<^J3H45
gNAcFXCAVE<>-J<g@XCc[[/XQ;Z^dOFS1MZQ-UIcWLU45FT<M9I7F+CbDP)\/YO\
I#XRAYa862C:YEc?(&2IMW+VdSCHX^L0SS=.+eWc);HA2MAN\-N3II5f]>a\KIZ-
.F[<2HHM1BdKE:Mc_L.D-)cHf;ZF8]T-]:[0gKBGS3Wf?YV+?ZLM4R^c2>)^=3=+
bL9N-Uf\W;JJXE=]/7L&^2H8gMKR1Oe^8#4FV,K\/6S(K5@N,c@?Z4dY2aRJXFOL
94/X1c=7VSJVIVbTR^3Wdb2W\8=M;RNa?7BP_\GVIX@aKZTHL?Y)&_\6_UbLEI1c
e<<>?2^\]Q+eDE>UNSCa76)TMKGSg1-7g#WeD>?\/Ge0>8ET,1G>/9VD.B=UM2C6
\&6NSO=TJ<:L<DOMJS7fLD,TVJ)B>-?BA<;9(>g5N<E8\[+H09X\Kd?C=W5^ee5e
I.]&MVK@A0c0)\P,IMSC[;V)6/O@I]bKRa/?&Hc_e)O;WAd3J-]1.G#[gSBVR+B&
fL^J4G.ZgAaS7gU=H&25=L<)e>R66-IRMES)OB.>=>eQZ+FS+TUcK2F.5/]]CX^G
PL<8FWVdF9W,0DGW@QSR&=B-O5#cJfbaOUWO6>9PCZ6/dH49WC_0(7(JSF0eIegA
3]RU(2AU/?7DCG@QY\b4)RC)@JR)fe@cfZ/U0J]2KGJ-@&6=[<gV8M1.K5DT8f\f
=bB=+W5>CP+^A[Q#6Y/I>37ME,P(_K_NFKd:EaNV=cY<1O&?#T1+N4I/LX9IBVKI
6-X&XRWY7AP,UA+B.RRC4/+2IUg(JCTbg>C69++I@5G)JPN?HA]HUPLcL]Mc[&#R
1660ZP&),KcE1WF+/Y#-OYIXBGGYI6V]c2Vf)42:6)Z,HXfI9:^6=dTO<@77L+2a
\HWeP]Kf00W4)fC^KT#G[CGS;Z9c<ObWeVU_Q3fKV\L1=RLMacKRUE;d\?:VJ5Q)
U2)GFK47e0=VP-)ZLg^WPMMS5]FP@COOb/C(CQK)1BBYSI<:P@YY(@6)gX&ZIE?J
AEdY)c@-99IJ:-]K?fIQ]K:TeX[VG:2-fM(O:,OB;.#f#/1W2?0eWN<_M;-F0CFN
#3_?<.V0QJ76@B)#VICOUXRG);52;Q^F0fC;696OZKMd3N2O@dX1]0d.?0@,TKO=
0O_>Gb^[NEf>2GgCHe&6bDR8g/IS7;(IPge44P#T6+?CI>B5#2R]Q;SEg]N=&.(K
=HIW_@(^e<?;7]MW/dCCK_PJC&eC[]<JQH#UB>:PNFB&<P0-@eLf3GI:D:aI7e=-
[^a3&gBUWXVJ;P9NY>;+)bbIDV(5SUM+118J#gA@9+]9)=V6OXA[G6;B/0JETcL1
eL;g5G^SU,K,7fVP&>Nc4_NN2_FQ(0R7_2[8.Q6VK.?R;O;:a#H:T2M]6H/V_7ND
3&&L@V=I/RYcP>=cZB(LMB12ADY()M?GV(FbDF.J/ZBMbF[5a45_,I@N]?_1[7DE
f#_0a;SICCY=gMQ08([?ZM<]L<,U[9&B+b=:T<RK9Q>g,&&>-,XLSgKJKf<]\+<L
f.b3VO:=3b68f_0Mc.K<62>ZJJJQ\_]2U3ZTR6e(AMWZ?6#?_-_0^cQ0f6a60KNI
.-81eX=UfaK@3O(J:e)G0[dgU1>9:b_K249f5;;D[M/((I\SQSYA&SO1;P,TF]eK
0dY8b;WC^;</:5#F[6aXeAb9HB@>]@2/>>G(a[R4APZR^#+B8ebVg&[SND=6d-]0
(/G=7(4V7Z,(VB,S<2AX>g7Yb1JU_D1:BZ]CGVa??M8V&R&#HYW,VO]=/K?Sa:0_
1:T4_89SI^C,g4,C#R7CR3-3Z937)\&[QSd[-I(_.J&852FZR=PQ,Qc>[2W]MH_G
:1,bea15/A5=_X9WZ,38N27R;#bG73(+8[X89;9M@-K:V-c:CN,b+7A&W>N42)?K
TJF+fSRHd,V70I59K6[R,:KBc#[+c-ReXA6:3ecSf3fDZ8J0JL6O>#9^(=<3:_]0
Q8H-b<)@E,<@WFH8a;O/5U3E>0Ze(-YFUDU0UM+H=G]_</W,[5:[SEf4F^08#SVG
W\>.SPI\GUF?P\]fV[=1T.7S<#TCHKUE2/cFM7dMO<Jb3a^7a1IdS7<VJ/C^/5VP
OgHWBg=>7<eU#aaVWUV[?<MYZ[eUKRf;^)(1WA=;>^J)[d(J.YfeF5V&?#VTDL1c
5bTHY_QA\HNV9AYbN#;ePS?5eEXM1(J=Gb4L7:?LI+d&9+;Z1QNF^DEX^)cDS-RW
+ENaCB8V1e\,eUP@/CC<B:=4OKGQ,Z(DGD5(?4+U3#Yg\_WPJ:eS.?J;,>>?1Z1P
PFGT7=H)I1?WDe0,2<]INR2:(:9R9WYDf(NK>CP66HQP[+=R9_</8D\V9<?JRBT/
@K=<O4),0SWe/6EeC]SG&UQ=E^>&DE]TbCf[A-LeBER:37DV/FQR(VeNK^3T=HL4
BW.+/A^\5\@WV;:TcBC]F>?S3L=RE8gTcdRYHd?HY)[-/6S>W6&bbcfUD-U@gKX9
Z,V]RKO&JfcJ<-:bHX?09[MSB6PIfa^;:^5[;F7(1=BS_GISXI>ZF12ee8?dWA?V
.[-Z.A(L-C=PgV[T^?1Y^86)0^DOM21\D_<F[;<#;9:F:ZYNF??\#a<O?73,CZU,
B1_;+d2LS.d+bS)\=D5_CNL5EHJ841_K_[?a[0FgVaX#f\W8-Fe.,Ca8NSP+^RT[
GC>-ZEX1=eQ9O\OOK6VKc]QKeZNWE^ZfY:=5c,2-A443;T#@=b7OF7O[eBe??2:W
E^T?GQNV,Pca:IB;>5:0V4Lc#?_FIQOfC?JbfBg0.I?YfLgZV#\b+DSSVOff@G(Z
2RED:^Gab&(.,&5Y6QIXPYZcgXc1VJU#GE]UP3gD;YRLP6KCUGS7c\e>LY#8XQ]7
03f9&00Y][bIT^4:#C39YU+OPbP?@QX5YRc=1F+(5Ib]<&N]gR?K:AWGg#,9UJ;T
\c?.=0EWC[C&KH.D5aGG9UB)((Q.@eK6@3+b[60?ADJHR+77>N&W3#MJS)KJ95HP
_]R+L;,TW\Vg)Z=\=S,Y.#5a50#\I5c43:U&WaQ]P&DCbY>E</OK</Y.eV\3gNM@
E)H1,S-,4B^\6ED_\:1Oc=FcC/8?Y>63Q#Q@C@7Db\7c/?\ZDZLDL,cY&C\CABN9
4J:[6FfR[-,#1gW(8c)KEC#b6<8cXVdKH]U(238d@X/9&g^4@7VfD+D8(<QF9R9&
P6E2P=U>TVF(^+-d=TUf5))AV_M4:7/+Bg54eRM^Wd,(=QcK;;<a\#5cb\fDT>[-
IcQ<_\W0Keg8LFN6-+9=S@SZCPHXYcJAfJ1;]2G]8)?DLPT7:dAdA.(AB-_QN4>H
+TU)eSY+&eE[I\1bG\II?a&5YM)W)2:R?S6cDdg20\Y4M>cJ;)J6()EELF#[]\<^
=COKeSR6^+;=5f]DQ3X21:cGRK@?K1^G04(C8ZgD;T&&TSa#O@[E5:4S2W]/.fT6
[)&e#JG2bU3@6_Z11cUF+3<L-66BE,AFKU6RYP8QEd9g4TbN+NBT@RPP(bI5ER.L
fJ2).FJU=0(RQ;0,bd7QQJB#8c\3Hf+1HSBd@HA1X.WF0<>RJ\Oa]JP?)?5K_eXG
J1L/gR8(-^f1Z^K(4U2G6\G1-+G8+Y.e1IR.^HEaH:f-GQ?JO),a3Mdb_<=,472a
,gC^B2?VZDOIBc2Z-ecEX+A?VQf6b&g>[gW<<5gP:f?4@AN0Pfd_.[2_Nd1B=78K
P;N3/^YN-^)1P_,WXEYAbH3&>f#G;d?0ORb<,<MeY6@7SE&41?//TPD\f_8A4gQe
(G4ET8bW8ONe8\SEFGG9RW)^7D>@JA9eL)SH?L7G3OTX8UP@34(G^+A^1+1V7,FE
W\MS+(09^LDR_ZN)Q:ZZUbQN96K,&D&7e+.Tf+XLB^/?L#gJH(.&TU>=/#M4aK&\
d7fVDeUA,)&)N_e(?R&ZZeLIL648^/f>_QLHgM9Xf&JG2fDLF;LJB4cgFA3&FNQF
fL7FFF]Ob3C,D&Hd_=[KP#S)WT\?+C6e((LQ=GI[WB\PW1e#\G/(aJ^G]QR1UPLU
Q_gcN:3b>N68O8_AAB1QJ>cO,CZDfV,,N\VR@SH.M)Ta@^0FY>bA@fZLRZ>SLafb
1>3(\^C?H:7U&)).;LTb=D95E^-cI0bO(UY\?)P-V21g(?#[RG7]T2PaRGa#f]:f
PP0AbSDT\9;PLb/YF>(&Y5Q7Cg,[aa-C=e[L4+CB@-F6RN@c4CD2b]16>-]NP4F=
?)g?gb7Q;Q+)=16]EZ/Dg1)]05T(g-@(F=07?cF2LV.KS7RK&.<#M@:-P]QXRGF_
C:31_6,JD)FJD5ZQF;6D4?RaL0bC=[5V[S9H\57?e^PaL75/>XM_)AW2H-SB[X<L
YQHWOF3\T]^>0:BC;;d&XWFNcX1CXb-34FW0XbK[RL]NW2<(g&E[fQZZNZ_0L=2T
2GgNPW,CH3DbRf\V1L@\7X/8\6dB+DJ=gL<>S\O_-CJAHE,DY[#DZeUH=C(eb4#R
>M1V?;&HBM,P,=OCJP,e<bfQgLX((Fg)fQL1Kd\^:GAdP6Y]1e:(_\VcVI;A\a]/
(f@S/KL<0@FAZM9+FWe>BTL_A)>:a+]R?.3(C;T2PN:QgdH,BcPYBCe3&3YWL?,Q
2O?/GJ/[e\9ODOGcTP5TSCP,R;SF7:=P=eaTPWC^G0(XSc=17L)eUe\VR)-V@-QI
@#O@Z01+[6>Uf@H5W_:QBGX61O>RW\c5^c6LAe]45]=a(;7B3GLQC/dEaDE2SITc
UHLG7\Qd254.E(MS1?6R],2Ya<@=[gGeJMR?>]=cMP5Wc@RH9[dG_06=N^CIUS.O
&5PIN-Z+MYZYOUI/eDNEF/A<H,@RLM9?9#SHB&:19I@)XV].,_<DI^0J.K:/:K+A
+SME6=B0HSG?(U<BJ&7JROC@.G_Q,SREDYP3<ARZ2M\eI]dBGE5#R4SG2;>S<A1U
N]VDd\=K@)g4:2U4UX\?.H/9aOac>15\/a(_H7A<2P;6,E+@#22Z7:+Z<KBaCXJf
U=EQ6H,V6=e9dY5/g_?+-5HI]GJPTCfB+KQN6a;\WFbJ9:PG[bJJN0KeP0L4-S>H
1)C\6(#aQPFH11:abATJXXdVf>Ve5.E@.Keb+e8:g3(+^@d;[6?0>,,B/H7A2GQ2
NK+G8PCRL4Z]dS58+@JW1===a;N81PaaH=17CbJTMa6[&B225SSMUUD-U,KV@?aV
1@O>T^#UC5>QcV7>?Q<=MQ)F6^HW\Ce<.42;CNbJ05N<T^N9?R\(/4,@G&gRS/Be
M4cda1U:PF)\?ZVNF^78:(CX6K83>D1>W3F>;&.fL4gfL,O97)JH(d\=UGB^dIKH
657?7A&SM@UgC8YV&OCOJb3.AV^V=D;G#UgD5/UEN^-?_;B84OP(+G+VA\d#X2P0
f08;YWV=f(Sfb&-,?XB(.72_eLdOT&Z23JJ3-:LdF+[dK,\3NWL9,?G:I49^+e](
)>->5OdMO1#;RE1]W-M/@2WA>8:J4He=[35,4_FNNW3V9]gC&YbZKGPWE3?gV=LK
+YUU(B)(fR\@;\;Q/3M=C\MG)FG0#XI\07A@AP[_:@+/B>IP790f3a2fc.7.SI+0
R&-B9@&Q9EP+eRGGK+1La^@KP7BB?Y83.EV\Q+Jc38-cKS]DLOW?MO;+Z+27#Vd&
>LSNS.WFY+8bBVHY(Y&RUVH\5[>dQBLWY\AI2Z9g,_7UT>3-L.;<QT^CZH?K<-1V
e17::38>DFbP#UHU3=S0B30<]d.9ML[<c7f5<f8=Y-;;(#<F.4F#A<P-/9Zd0:JW
@eJ(RU+H?5ZA0>P6&YV1RB(g@AM9Y=I#]L;-GA9fX8S@T^55PSC?(,\C@=R=(:NH
-1Q-XHN2G9Dc<;PJT#VE=)G_bAaGFN<7DYXRMPgTO:[5^R&FfP)CHR(bHeHf6NLC
8M1WIXQCbV+A=AF2X7d[ZIb0E,?PKV]2eL)/U-(@WAd9[3Hg.(;TCJ:(Q])>a.6/
62bHU)a,2+<#7;R;4YH+;5+G&EGKF5PMRR3Y3^e\KD;c&a4e#M=&TCec;ge4Q?U1
1;#J+1V^<Mb8Z_HI]6RNA+W=0;U(2WOf2U44L4\dd2ZSXZM4GP)d(Wb7K=Y.@=\F
bJH^B&YIJM^3(-S]N+)4^;09cRKXU]15f1H@G;9]Jf,DD>9M0<+dc?7R+7A&:=D>
):<bb,(<M>9#73AW@SZPIf16?gP;7]QeS&:RYX-(7KRS;IIc666^#[;M27QfR6R>
Q0AD:F\T)>ZQZ_4\OK:+Z_NISf0-4b/1\YSP@MX>DeW,3J4S\f[fL[dU\d:<eT/e
/3)M)A83VGH7:)-_ad8)Ye<,();^_XIUg4/<U\U/D,aOZ9R](30QRIcQ;8Y@g#(\
S-S(A(R;,?<ZK1aNb9f^:8(#9>=J6_f\0;/4(7>]d5]OXW@_R,;7ZP<5N-C3@[#=
.^9[,#8e0MS.aJ8BS+O^[IQ6YYIEgbJHd.9Y)5CgL@ca<FLb<8SHY5,_.(-^9e_b
Yf-K60-<adPc@O.)1AN_gV6-.[7<Z57EX;)Rb>0-#@KZ=H\BAH&U]0]9>XT\=</O
X@4H_ZL#/&0R+>K2E(;+OdW:R#4M@U3+g4D<:G9G>6].[M#U?;KPPE4;Q3:c<+8d
MXIGc.A/Z+SQJ[(bQ:_9,Z<S0/Gd,AZ16f>b=,C6NPfV5>#gb0#?JVg=3I[cIX48
\\Qd+cWJcD#+8D+04@La&C=g/4=RRSBWA(A8dSGM0Z]/dOXQ0;RALFBHbN,((^Hf
;D(X1C#-W)^b8)KQ1^3KHg#?G3cN&B(=U>MF5LBI@cO8(_4/Ag[7C2G2&XLIgBTY
f8DHC^BC?V/CZQ<^Z5a/@(N&Z=]0(8F>OeMNRTN^::VI1]=9GJ>fc-(^H+#:8LQO
_,I6<2/7>806Og](1e7/.^^8>/K&;8[GVZ1d_53GV^>I;dE\FBW<BR+E.L.>@R7=
2N&NHR#bB/J[g+X=?e3XH9/Ibe6E-X8AFNZcU\\,ZA_E&ZDLXac1V9FALAFUFE_E
Y,#>33BO,A[ce(@ZV83L3PO&3:A+:gK9ARR3P@ZNE3C\(+9E98/^WF8J.N_F?Z:I
/-@JB8aOLO@1^TH=1MNb)QW2-X&I._1HKNHGBEE)c6f&^89S[@1eME6[LQNaHcN[
\K3T0<S.6=V4K4B8W8W35:5<=9^-:Y:^NdYR:O<[/G0I<J(+eXVM=5Z6;]WCD6\6
7a_B0AR,QFXGKXXge3X+D/?@0JUI9A?>aF<aK0@9M\\MBY0Q5RcH;Va.,?I2Z5_[
D^W;dV#bL)6-:W?ZgH)?dY+6FKLa5Q_X7Zg<cV_]XV#RB/.<0J,f5eT5,,MEfe_U
BWV#W-@-2,3_OK7AKTHSS2@B0QX5T-[eeM1_.M-4(QSHK48@\>f^U5gCL?d<g\NG
&>H8(K6CUgO;\(4ULf7:7LT5J<b\=IO(KY,Ped@Ub.D<_T0EWL(\fF0YB@<Q2b8D
J]SVD+Eg1PXBT,53&7>8S4A,-^d?U+)0VV#=7C<)JVW.Y<0(_^_@FG.@Q?Oe:<e/
UeD)H:V1U1-S\ddI,F8eAgP:[[cRBIKKU^a[V=18MAg\1U)\3;9c&abRW;H6O2ee
P4@2E^YM7f1H[VA0;U<+P@:Z;;>[8&@U7M\C__A2<SL3S@]e1961GO]#@C2WZ92f
<J);8VP;C#-->KM;6&0EAE0]eW]6[3-AL._Bf=2G9+#ZK(fF>AQH5/caEL/Ueb.&
\\aCHYQYNa,\=[<AFTQMHRPUN_d0WNLUMTgfO8Md\<(IV)&C9(64@KC/f(bQSIdH
M2\c\ZIQO)U-H0D_6R4b/Q4^D9\cM6ege^,Q[5\Ca(()I@I2Jeg\[cB(ODfVSe]2
PKT,>>3+:04f?f0.A].X/FZJcEFY]NG:a<6ce]ZD^gBXV&;<Y.eYR&@DIVT-HK5E
JdMGCf@aO6U=X7dAXdePQa1g:.PH]2/55KRdJ&CGdGJ_W.eYKS#YC&^c2DY;V[V2
Cged^_&I5Y]E],J^<>J(<JP6_,F\OUK,C(KK]TQ0L6cL[NXLf93b-69Gc5eYBLL4
B;gDPDZ1+OdfU/@\f6]/<V[;Bde\aY[P66NeW0IOB<SV1T@E-[NWXFJIb<OR0bNH
V)EO0)^BII+>\DX[O2)2HZKXK6BbOVPIY0b.=55H5.P=YP_B4^&P?CK[#7H_aQKG
/2D2bPV@O>@^?H8FeK5f@9J)9&?<2S.GOafd^2aER^.b>Gf\g9Ec]VAZ&A7S^OLB
-H3f-@/c<W?5ca[/dO3OWe,(D;-RSa><0-/J=1^6cUZ^N>HNWS)D0ZG&,BDS1aL-
VS8:DX+#g,6.P35OVfVaX_\I#;#<3fXC)3UG:)2&DfYI)+;/;TH3P/GK(>cAKINL
LZ7UNJHE^STO\8V_fQDH9#3]8]@cIZZO3,e]3H-8aCM))/SBG_PFB(dZ1&Na?4N=
SJ[?-c0Aa4GPH2LY:]OccDE8E]CeE&N-R<_A+^8,M,;),1@=3UBGN[WIUZ4Sg;N\
,@B]eZc,Fb&.9egLM8#GV9.P>-9U-;T+Xe[;UWV_N+Z(7K@->&J6OaI#I-]\IbHS
OT4U_EINHe@-1d7@d?0c7fg>BPGJ]-0dXfMJOK2\HU^d2Nf@/FRL&E_ee/2e^Ucf
\BQ&ID_<2#3BGeS4ARML=&CV(MQ4B3B(D/:W&.VCG@Z9W>4EbO,B:CeK(@c3^0(W
6Cg(MDUIg#IN^J.SP<D5aK<4P@,Y+27G<VcWK8H.3]Z+e?NWc,&>cB7Yc<^92.:T
W<M7eV:a<FUP+dS+2F9ST^J60208eI(5BCL;YQ4f@5f5R@1#_Ja#:[XWDHD)HZWA
ZBVO]Oe688X,RZ::+FAQ)/8+f=NAWC+O,[FIMe2_O2:YJEUaMHaNRL9:W9>D.VU:
9G&1;.B[:]a(J/E?c3:P9ZLLM)>6fTcI+/8+ScY;.7Ig_S&Bf]2^Q0Oa8/>2eEK+
2Z:cR0Q3-#DTCBG?D>4gW3CG4UAX;HHYO0&2WALIZT/:LP@\/CRUE4]cNHLTL#\\
A-<D20,aI&G_V+c1>RK&ae6b(KJY3a7C/d]\49XMC)Vaa]1L&^_X7bF8LITe8[8W
1_8<?P&]SY3\T7eMRQ#7DL,4d>S?VS)^7VSXX(64W:<9;HU5Y,(CJ&8Z^96b]EbL
OT(,CcW2NaOS&Q0;.]+Na7<G_TI)5N9Q#EQNeP8QQCWE?F<cd=RXTN-B9FV7\LFI
.,54HBI2e-a/&:&P_PZeM(W]/;I6D\)C/7_cO)#;UJg)D7DR:5=665eRb4<+=VZO
NV+8UQJ:UD>21X>-aRA7JY4GfO2P:ZZ#e<Z=dgAWC0g4P]EGMR9BcQUd\7AN?I^1
1RJ8#5V9OC:05]/81TT__?IPV]-T/f9[S/QaVb2\7Q?3QcH(9VT,,(B#LEY+\Q+C
23SJJOZSV#_SZe/@MM_PZG]Wbf;gI0(f<\,_)DETdb#Q>ZU+)E?e_LM@O^89CRTR
T@9E<.983),JZ2/N3@U@92F0.IW5:cM8N04g=:,>7YTeC.D0#f5AAf#K]>4/17W:
D8fd9F5TEY(1\))W@Bc)<G]2WGK^@]<>@.<W065KL5J+ZP)MbK_UK[Q;MFO0Y3:e
2HJcGYOHCXOQLc/L>3N@=PMQ9g_eD<F5T#8b+cgZ;PB>DVMB5[](Z,f/7FK&IU,X
0G@0S\VB,_KX\N=K/MKV,:)XPcUXcQXaXTU:[@=5+-H&S<B_49KQDBfA6G?W+[=X
?4@.g\V)?5>;eA0S)M\f\b>262^,B&HBNLc]:f:-4@TV^C<>&YZdgANM@\(fcJ1_
VRLHc[3]DH824b,DM/P_AcZ5<J[BK68^_aGYB3L19@+geC7Y28()AbWVU.FdIVBR
bf#d>JCZ8T@\LaW/OSfc6EOKf^2JQ03aa]/;[(0UObU4M0PR.fBGgI9=4-CRcgI9
B(E)S/C^IE8U7a:<X)DgMS(]gf+^B@(S<82<3/)314H_CFVae+]WQ1-,NCQ&eeHW
KMRI?<Z0E4@YgQEIX#Hf7eT6LN:U2/FAQV+?e+)@_Y8>_5N2RO-S0^<R9:EBF;?X
(bH3WQ-@]5G8P7QaC3d+GU(Q&f&TEWb8)^/+5A;0=3:6((TKQ8b)ZQ)9<>4IA<)R
PAYgV:XFBg?S6(YL+cF\I1G1VOf?Q;T5\VQO>UT+1;6]e.(/,Ig<I]]#T9bCH+T.
X:5c/-0g1[1KfZ_H\;)WFRcf?9&68UU;a-^Cbc.aQ4S.d8FgH8>dMVN1M5DF@8>b
N_TNEc;>g9cMCRJ2TAH4.d\dC0O><3(XKG+b-aU7f.OYag<_bdLTNO8]3&Ufc>__
,HTL)1]=JCA=.4TMQCI(Z1JD)V4#Qf38RU_Me\F^fR^9[=GNP_/egJ7+dR2:F;L8
M^]GMKW-WTe]82fF&5g&K>f;\f=FEcKe.GU6VQUV(9NQE@c-18fX\fM?RG?K2A/9
ML[QZ6V-AF>#6/TM,)O3;4=T\4bH^]6AUMJCc(FPD<BM\N0Y#?J=c#[(:f&A7BR6
&#&HRKXeGBJT?3O&LcO;Q22A(,BdN-b.[dOC[2\feV@P1\eAc_&T;51AJNJ<Q1.Z
=)&LI7P8J@,V/_,N1<?.gG]#VOM3b@8@/RVL6RD.12fSc.KWaf1JFJKN7I))g)IO
4eYWPCEE/MT&@>Z89P_fP3gB-\d\d#,-QG,EM8MN=KE/1dB>MJGTM_/SN:[6VQ\Y
:1>_\8>/;X]Taf4XdEQ:@4HS;=?B,OER]I:dZ0&Y07)9-/4XFaWT<^cHc-?B?T4:
OdSEbWD5X0(8[F@(>(7(77FQHcLT9RNK#-]^FP++bCO/K6d.dJLR^18f/dD&,a0M
,BfJHB+[I[7&d#Z<&SHT<feE+bOX\(A\LQeO,UC@\Rbc=)BCNZN.R?-81G?d=g_d
F#a_IFAe?.+f#,Xgg&fBK0Qg_XD?I=cV0W,L:4P]\[TH-RFQ]a^PFcJ&a/aFg2MG
1+;=P,gE;^-cET7.(Z-]af:ABK?YJU7^T0O2-Yc.O<^QRG][;<<]T82N=C@T.@FX
MfL5<V+:T(9Q<918:=Sc\@D.OV[T&@K1&EP7_=L#+T8#49eLX?/.@G.XfJ,C#[<+
#\gL>)dX]BD,VV:IDRM3?QMB6IMB?ac(&&=;<Z10F=85bUBY/WXIQOPUX,T7988X
Kd>20/WYSUeO&=U=AGNS?0XTaEQ0\P+g&=Xc>B@[_#ID<2&<e]+S,dMCWF>_9H9F
-&CED]>8;L/]]T3a[8_RI;1ga.(7^d&OY#KZOO^ec]XO^,-[M,KNC\D6C^?VO[ZS
COS@Q3)=NDP:8K)C1T/7M;-SVWVgI<?HB@d+KU-K=6Ad7-Re9^VRKU05C/+Tg5P[
5Tc;6/RB.[M:9/I(MU:CZg?cL5NAD]&OER@g\D2_NGS^I\QC.Od;P99,3^J/e&O&
g5UXV-.H5c+U.T5)+c.(8H0cTKe>V4_fd#Qc<;IV72LT<228<d4A8SWdf=#GJa&I
R9D+TcTUY9&(&R:gc/W7eW1EPbZf/8+.R9[a3R7B[IX>DJ.f[^7)1f?1[+dPbeA1
6VXLHEfE5]1V+;;B<B0c3[>S-9JQI/8]7\6S3NWLSCXWJI22P-Z_8e4ME0R#Meb+
E#4)>CXH&=&<AQ=+5)B<0^C,:91:gI#74._Q3LB<V76&5BFe;[Z&&dAQNaT8_B3#
5S4;TVE2aWI5O,cHB4.OW0@S=,IXNM?[C8F@)D8YGdH+ZYbfY@]M#X>-1O8gHTIA
D<5;0_^S(78Z0A(fL_g-3fZTKE>,>IU1dCSOOM=LXZ5A4?;T2OGf_g1E&4d5TSLZ
R?<_X\-LL]=a;Yd(]<ZO1=&P\gO9>U?LVDKW2@eXW2?2&5G22d[6#B)S_PD\U2R3
>G&g57^N^OUZ,LBU<)bQ(2;/.eg3R9ZY:9B&W=d,=[cg#W(XW>7V:YL>C00e,K#a
?(^[Y>5P=V4N4P>U4HJ:TbH2?]f\5O^NROP](PP\.>MOS.LOETJ5MCJC2<M&8+(U
:^d)N)26-GdAZ+Q/<1<GR-8UO>#Ic@-AgD@.OG[^#R;1<.c;3R(=fM#(KB=?MRV-
EJPT>UY&S)92<4ALV.?XY.]8FbQMC-c-dB^bS+NX5L4WaFeR-/JHB@TQW7^S77E>
Y9HP@@RcS?)T:IM0.43N+8b)e]Of[424U1W3_)1O:VM3WbJE\64V4(-Ree=4S;-[
CB;[Q(KcE=-,1b)WU,Q)=^I^NKD0(E#QZAKH;,ec^SC2d]IU5O)dfID[6Q1Kc&^1
Y26ZH]S6GE[^-V6=NbI(TM8#c&&?&S.cWJ8gY82P5CP=FNEK-(Hce:4+GS8/dR.(
NGdJN,SI@]F(-W.A1VFec+eIDN:+<R3;69ZWaSdH5d-&A5^<<G]Ke.]/5\0S3-a-
9RB;?c>)1B6CFG3RTZI#CUI.9&1;:?-AKMf<Aa3)Fa7[e]f33]OS_(#JQF0SWM[/
I-HV@]8#E_a4(.LJc1?TWOU8bOH2#&5];N#(e-I8U@WLFfM18,fV+dQ<<\U;Qe0C
[J;aM]9L8PeQHVd\5dK=OHB2eXJ/K^@>WSEf6b92Q[0N83a;<XH/c><SBNNNXFQ:
APR-b]^87:PR5?S_)NAU>[[5G8P@NA/0Ng;-M/^g8GVF?e2VF1L)K(&2W<#[?58W
R5W?V<JRX8>?@4IR_:Ge;;Wd8(O#/47[._a)5=1H;+Q_)RW481V>BZOJgdOI)/F@
f@bC?bA#(&)12g?&Je9J063?@5MR0-)=<(W5Wa=JZ/Q-\M09NNb1G,MdeE@P#0A2
gDA]C^EegX,)=XJ8><?PT--QR__<GH0+e+X.SXKKM,c]Ye3;#b?UHS;K6f[HI>8W
84Y7<)BH&.3V1R8,Q9&]_cbD:Dbb7FLE=SNcVG.Ce7_2:[=PM7D4,E]^P7;_d?^,
GW6SP]c=?<R6X1=@;\NDCB)MVgbQXWFDK)TTTOMV)[fB#VKO_O:YG9C=S>?1KZ)^
9-\H\//6_3da0E1UdKI[@H//=U;M1M\F>Q40,e6]-H>edZ7Z?]V]]NKA9JK[<c25
PY;^.[NcC?W>NdY\ZQgFZUUP-O3G#[e\F1(#+g/]1#P7)73fKY3e8P>KB&O&;M06
E:d5R](^?BA/M2HQ-J<T^:?+)YH]FZ:,DR:TIGO^]8?>Q47O]>9+KKZ3Nf6C&Ud#
;VMT[4fTA-27<@YH57.g&&V<BR,:UH;:22dDU,#3.Vf]GE9D1PK_g.KHb7=f>XB>
<8\:HM3GIP#JQCISQ^;P>@:KY.FNc&J2R7,A-R6ZPbgO9+<<7S49.0PXW4=Wg9-1
,P]1b7DPEXOW7=@XN\L#.bMHCC@b/Mc13c<ASG^CFU,[;AYX3g^ZBR:3DL44ae_I
6ZeXH&eMK<N)+_Z=[D4]C;A9(E9g9cgd9[^H3\F^(_e0P^>WTOaE7)8:Q2N:O/D^
JF3TO;[#;NEZR-EWQ0#[1.I7]7&0\N]YS5PbK60CW2RcF@@QdRVQ]\[4UG+(Lae:
25?O&eSY5RY;9;aM=-HXZ++.<bJOFN1<JKQ>PL,b)6+<:7SK\A<VNK@AW-=1.1LE
d30f6@X)8.I/XKDb9Q8E^Q1_gS7]G0WWOb=0U+5f]#CH3g10bD-01(b^SHMTN+OM
/83BAG<&.-].Jf4+-LL?VgX@NOLPF;1f<XFAINDc5BdRE\]JM6a&OYBA5#H(IYP3
fXPRYY:W,K4]<J0D8NRB?IQe^d69?Q@Z7BgU>?bU1IgRWAHON[&46#@P25^4bcIR
.Z+E[MCTJDV.RQR;D<c5FBRKGHY]EVYP=5(2@5E(803;06g\JMAER^ecCTF+(4XM
<UR/&7+_c@?TYbddMSd?V3).4MFR@G1dB3d,R2:\?Y]ITWacBg]._AJ(]WTKAY&a
HfPg7Z+N.d(PdV-VKPRR6\QQde=48?)CZC<CE6&5K=]0c_/aHc]3P<LJNETYJ_GE
cH=47RAKD<\NFD8&8#LF1N43.,GZH:8FD\.L&MEPPd[,3=TFYAQ4\#OF,[V>@1/W
P9X)&V_YMDT5)ZCB\N1;CP+:V4;UTV#-f/a)S5W5L3G^dGX?dFRFM,<MSL;+6dVD
f=9Q8&AYW_I2D491M4BGIa]<52aJHbe_QKQG2H_V2gM/:HR]D9&W(8S)[^_S76D]
;f+Jf.2dLFMYCR/(/)D80539PS+5M0B3?X.,,_Z3XCc&=(+PfA,b\P@UbG6S1<_>
<T6d&D+@T\4QL-=1/&4F=4(H&:)S989_eC(DCJ]MPS8?W^.]]Y6T0C_\R)G371Bc
PZ6g_)2C,.e)42[c(8BN=]?U(HK]2a+5GLNb<d_&DI@G,OL9Ue;35RA0)cXRFG#I
WTA_8cA)8@g;L^TcIS+XJ)M_)+I404[FZJLfTQL40\V];@B36+Z:[MR99#+N(U@d
[7)GW@<C>b?I)9>:)\G_)-46QINXEG/D6JE+XYY\:OJ8I.RTO?Oe:O&#)ScX[(;T
9NS/21:b,QgVY\d8@J4aR7PUgTXXHdHHEDUX]-8D?ZbCU,=^G=VU/-G[8MGdL18a
_b5D&,a^18N2M2#P_,NXf-FFC>D7QJBD\>AAM]^..WS<K;YCOV;NDg=5Y?88PZBa
5;KeP]_e@9LT7&ZDY/IK>2SN[4QMbW^J.FV]Vc0;Y^.T_(J?2a]0SJ+,4&R\)cGd
c7<@a_-WC\V5)7YM_3^+C<f.H@]B=a(42P>56F]]_ebZfV:W)(gaK#5JFeDG;B@?
C6=)?dLM70gaG]R,P.d25(>W-W:8VcA^WYN5#Yd8YdT:LFEE^)QB_YX+LA>RBZ2X
\+4RQd6)L+aa,:ZcaK_62[BcFW@ecH21O3_AM83UQ/@+QaH9SDM\3[/(Z8S3UV+)
^:</LORO>ZOXA?6F]OBF^Xeb_g3C<FEF6\/C9D#B)9,Q;5YJ5dD[&/CB]\5JFc>7
(E@^Y&G;YES\4,Z5)#S(eR2b>@D]&3^eJU_T@V4aAPYd]dOUZc&a2(4cOC7>0.Q;
5FXY5Tc;:/TJOdXBO6e8QHJM\]^7c]WYT:_]+-/NEN/=ZLe_Ic4>&g\_R[=<SgUL
PO4W7<,DP6b[2=E5f)S&cWLe\ccIO03FEeK81R7XM]\dPR/ME&SRG#XW218L##2F
CdHJ_#JXV9eP0HY71;\N@OF2d-#@Ga[QY_0WA71]8I0DM#aWa0M<8&(NFHSW)E(5
WB/Vd4AdLC\?ZAgGM,<34DbD#?1F9<^P6XE9/3Fce=d_CYeM:aXO&M3,FKa&fQT-
=8f]<Bd94b34_8OQCYER67?GFdMULF476\c:bSSHX)fV;P?RZ4V.C>ZDR#Aaa5\)
RcD(S?4:-^]1g^b>IAaHf=@<1G+[OK=@fgaLff35#.#F5DJ&G8P+>?R<49PG+\Qe
[RROLD;g?(3LOIFI^Q4T;-(,dQAHTdO-^I;G7M4JH,Uc&:EO4b8&I30SfdK0[&S-
#fY^AKd(7V&Qf_Kbe+4X=]a?TDVQX[^<6f1Tc9U2TNG[eYPMIQ?@[)IETQ8\:>/P
@ON&FcRIBKU-7R#O;(T;gA])H;H)\]B\E6_:0,C5PeRX(-W<6XS-Va1daQ=0?4J>
+PJE[=>([5,ge,9WfVe+c:J[&VZ5+JdA#b3F^?N=g=WR;^Ka>\+UR@74UZ[_?HF8
:)X1#L-[BYA&COR_I&D;TE.cOg4OQ1IXG/2;ORUX&<F=f&C15BX1eRC+N6^N5VG)
5G/OAPPEQCAW];[IL<MKK-9bP2KI,f18PMOZV5A]e3gCSOPY\D2^e#Ye67.8+Xb/
/31?e/a[?8N9P<4OY_^2#&fcJD9R+?OG=-<T^35^JQVHYaUKM4f7C:RPXI+B9]K&
I9dHJ?<_(K]OPQVS#5P-X]N??]>GODg]]:J9=EPEZPV1(<_/eZ;/KMHPB1=Y^):4
/),UN92\J&Y/6W<CZKS1D<E+,;F-L+b,=A\:dJ8PXc#Y:YDLI5J]?Ng;R(0J4D57
=9bI&J>J1MJ,2FL1a8SBZE843T:H=6Hg6(RSWCO\XA96G#G9_CFB\0+bHFeQdD:b
#YF2b,)Bd^4_#6_FN)a?cM27IQ9>=^g&bN6\OPQ\De,WCaZf4LBdXQVQEWQ(D_?@
B(_2:C]]f4Ag2)D[1F-71MZPTHb@+&_[MN2C?,XfW;32a-?W(WO<QE;QR,&E[&S_
VE<B80a0JIA\S-aN\720^G9JAc#Lb0Z8;>8>P531WA]Lb_IU@J0..Z-OE]MNDFEB
K?<5\7?D1S?A>U[5;K[&7QLFN)LU;0/7.>X6F2aYX4cSXF(eQbM@10&;>L]-=QX\
V<&_H;=NE_0&-OK#a+_b:<=_<5=[BJf?cAEc)XOZ&OSfNf2M_&0C^-:2L6>)Rf.#
Ha_IF/)(KYfeLcAOg-,08<U@Z]ELJb=H&025]^f3(FL<e/LIe)7)?)6X/b_a@E>Q
OR=R]VY5We:VNQ95G_BA;,b<aT0bKe@):a#XVfQ4X#(5NKG\<NdG?E\OOZT@:5]X
37S?74GFCb4)1TD?@CSTFad[MHZb\IRZ<Ia;-GSH1QJ@-W0CFXAORWd9U[#AO+H]
73P/b9N0JJe]0,8<XYaf&G_2?Sf1cFN?1#1ZQ_]Q#D)4>X6dYeQ3FR3@-]#8d,I?
K-.A-.;J3A#5ZaY6JgTP+JW2O2.[+:4A3/[8D)G,bcb7Q&.)bdJ,a@IU.E9O&=7B
=\:ZNA;NLC9XIV)?^G&V;\/O^7GYMWD.5gQETVC?:SL4eOCLD^57c8VS)[61GS-b
IbeA8U9P9)]VH]a]01U)(OENSFPGL?Q&D8RF,.+DVRNZF03P;]SN+:VdV8GY\Ce8
W[4J9a_U>DRfP+)M_eK_.SOC__M4SI0\#_AF+?QEXe((EEM4_HC3[=O5<fF5MRJb
V>8)a)dZ^8>ZFb0FB)6DX&]Yf;2]-,3+X,^D(cI5KGRa[2L(ZSLR#(BbaNBdgc7F
#D/QR>MZ#/@/>8U3(17gQO@0E0TDg+=gEgBQ;(SL3V..L-ga/?[a99KMA40@]@8R
9eMG&eW+/+A3FC@?(694#2S0cR/2101deB19c9:;bP1)5)f,-NAff.<c0C6#.fZ.
._<)A6?@T1&fGF8+N__Z]0BC6MM].D:)HKPG)WYOJ1c/M-+g#FMgO7R;Y-L4AJO?
H+fOHA/O92]>Z0#,GL^M3bgJ4(3SH^cA&g;NDgH6.WaUR,3P\?P<,_T=>:60AHB0
5L&1B7f<RY3;9S(fAXYU<f1a]IU0\gU+cE=Pb1_7:/&d()Ye<AB;d8e(5?e=VOYS
(2,8PH3^NFTNC,+W&-@bT;.Q1FG5AP\+#EPg\ZR-[g[@16?(CAP7?ISR-.:G&-a=
0(&f<GCGbWA06^&Z]HeB9EFLX8H1RI.4+86Y41(698b(05TdRU]Z\3:P)/[RfJgV
&;@DYGV1Fc3NDFPA9ADD3FO\?K<&FS8aN]OI_>1F1[?9/f#dMVOO0GI1BJ)TZ&Z6
28>+6Y37B;@0&I=^IQU0bc9;+YRM/2EF.N7?L6KVBH0>Zg]757L.94+EBZW-N++;
dU]bVOGJU329Z63#/:_NC[?ISI5(R:2&<I)8IZBY[0;f/Rc1d8Z+S&NMdX./I2NL
e3<EJ>M?<Xg_Fc[d_aVa#JN7(ZfT[&_&Y-#gfKb5Z6/?JV,0ZYd6AT+DNK:B#@Z+
_45[7U]3Z-Cac6FOW\TWV5Ub:1F>YdgeO6ANK0)/WI-f]40+Cg3R=18]H-agaA(e
K,Vg[d5#UI<BaW\_aPaAG=Yb<IYZO;WH5g#S[+W\Y(,:3YZW3[ZO&;3c5HTU<NQ\
8](US4a>M=PZYYQ:.0UX?TN#;WQYBM4g=&R2PNH6[4g2;S)Ge40b+)KQ]=\MRV@P
3f29,-d&@RE+Z)?fF3I^b&>BB1S9_2C#7Y>ZK;>1MNDWU.g@1]F_9J9FAAL5-OYJ
@@<9\>/KQcdXM=.#>@NXYg<;c_T0)fb\@_\LDU4JRb53V6:9XSDTaX;]@/PG<>U7
gF3dddVQD00f6gG+722&)VBObDb^T]Ra17-/b6-S?5=16+-Wa7^W_=_CB+VR&EXU
<)P8,]O9#ScgG-f#44E_H8-f:IF)fR?A,cB1W0e\VSBHF]I<gP1K_)<fNKcS:#HX
7MbJZRC+WbG7>#EIVOW>[#X==7[E.<8UF,BLM[1I3Lc<g(a&0g)7)MB:<;OfFX?=
\bMXO:];Ie.D@)B4KfPCLZ7TJA0@FE(G>4Z8F?K,@3)/INd50(b4:XD,Ed1VaI-3
MgB1QeJGXf,d=/P[gCMdWC+.EGL,d4RS9g74+^YX5,b@@AI\&S>M][X>-.>86dQV
&KGbb<-I74ZB);34[5D_#V<CgCEUB9e=W;D(-PJL^BbT>KJ_g;H;c;&d(A&S?07?
OH55X\ZBD81Me^M;PYN,5JX.4Pd^8e4QFWS##g.(;Af/;A1<.)[3)g2\^g8).;eH
de/Mg&<1E/#_/&]F\A<KNT=8.[Se.ZRU?XP&eb3TIP1b3K5:c80D:6-^]7c__a&I
:Y.PNVT#Y>-fW5#R=]BDQO#O[G:SO]4JE9=??#FZ(.EW4)A#8\V.>d(&78-+)WVU
Ugf2FdZCA?Z:_0+A+Og.3G3cUbIgEN(BQ9S2QBE04<200<b&(_G[IZf-<P?D?-b4
c]P6>-G2HZF\Ha-gCWH=XB_1f4f,^4OgfQ\Z2-a(^0ILPT#X&:(XX?Ma4)I&]INZ
]O,9RI6fc+2/35gHd-g<+R3G16B4+f#OK#)#E8cF_Z=<Da81DAK).OaS:/\4+?XJ
daZ?RQL:3eD&g-NTGdWHK0)C=JN]2VRJ@^#2W]6./WUbfeM=4]g4c#+N?dbV)bG=
e,ed:e)O,H=[MM40(#A6f^b?b&SQb)aAJ@<YD/Ec1gaaeQd,+.01C4[?Id=D3.?e
]:X7d#MBA^+^RD:SCb=@>a<-GaO/dHd]/:Jc?Af_KaXFW_:6W)dOY@39b?[18H]1
QF;+PKN3)g-&_K.908\T=&e16XP[,QfK/-e@cS@G>J0Hb]FL@fJ20BbFf2<6^]_f
QHFCD#SR@d.0:-]YGAT3J5.-E54aG8>H;;:?]4b3C\e,U(W<g4+\\-4H3T.8H@T>
RB6CO9C?S&W:0+)#9..7T5X-gMJR2]CeUS[65Y>2K5K]3OFWUb0;TeNG,BVXfgY=
+P?O2_HS<DR=I@+2O=(gHJ2OUeOSC;WX&NJc6><P=SD)A(7ILN:cK<C)X)=D/68U
acQ<eTKGV3NW3945;Z22^]cO^?R]T(?@f3.\).aO549#F^T[YRIYR+9c?&(d66Xb
0?4N-Cb:[g_6OXQY:O8bJI\@JM+AWb-4f8(TQbX0.1P1fA\?bW\<7Q6>\=AGTL?P
5X@EUCJ].,E8.+3X]]PRH;?,&U_(53J\LIa=f?aA(+J<W__X+Y9,5#3(P0/TMMQZ
fN8>;C)&8IO(X\]YcSZABM[;f/H_,&1)SFCFMAcA3?eXac.b[]-XK#.a(aG/+7NO
Y-bTeC9V2138?9bXg?dR0AKK0/I?-I,[YHY#G0[FVI<+J83O\_WN^I;#aRBTXeRB
D3WANKZdOFW6H(>VU4=UDA0MLDBJ1QRBL)=@@^Qb&Z8VXGfDO1F^H.#bFG#C40^9
YJ?9GOEOgCB7N#UW[8@=72]6B.<NRd3]c-@?S_cG]G>>1([ZBY)U?OZAKW+Ze\@6
ceCMR8L]S0VL^<D+P+5;PUKA,RZ,DeGGZWK_BP;D]?2==(F4?3TO-F=1@1:)4Hb9
&:GDW?S0;QQd8H&B1U@0f(B1G:R7egU6FS:/FL:cH376JR).4^TE(D9TdfFUN0:?
-W<b/HIe8g7=N7:I0b<>EeGU,-JJ;_f76L1dJBAS3>2)R2?e7B(KK06-_aLN7\D4
60VXH<Z+:2G;-6=GA1gc4_dB6;5=&PfTQ4?1YbcF+>b0XA5@EdNcZ\6AX6:&:LcJ
]>c#<eB0)]/9@_]CPYYa6?DAH,WY>#)EN>O@Y7>M3P\8\PB32CO6,K,U0eX]N97;
XVbX?Ic3^7<bCgEOLO+dC)8/P)MQ+IgD_<&P8aId24L7WJ-adBL6LSCHdEP=G?G?
=I7Vd>Cf:S\)Nd_1/]VQX]0d(@72g4@VXGCS[A6G]V_PNHK2#Z).bM.D4LA\]_G6
eV;ebC4^(^QbE@.=J<c##DS06g6eN#&gDdSGKfaVRb@W_&f9^44,.&Q(9CJfe3?^
DXe=VEQ-GA9933RcABaE+7FWO=C)9[A0c4YN4V2(A<170=,-GXGdNX9[6:0C5CfH
[_0gUc3]XVR_JXL(QQcI:SYa4E8];K9C50\YeL^:UMG:L8K/gSD6?D_-fPANb)T=R$
`endprotected
endmodule