/*
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NYCU Institute of Electronic
2024 Spring IC Design Laboratory 
Lab08: SystemVerilog Design and Verification 
File Name   : PATTERN_bridge.sv
Module Name : PATTERN_bridge
Release version : v1.0 (Release Date: Apr-2024)
Author : Jui-Huang Tsai (erictsai.ee12@nycu.edu.tw)
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
*/

`include "Usertype_BEV.sv"

program automatic PATTERN_bridge(input clk, INF.PATTERN_bridge inf);

`protected
>YDIN+g@L=?0e?D<3DdMC(VfB]IbX3c?bL:GD#0;)D)/CNgMLL_[-)d-@W?)f;?W
6CW0c7-6?fV=)9M(3CJUa.G/0)/WA9M?eMXgLH8<E-SZ;>Z>Ze+-U:5[80Fa&3S]
<XId.S;4#./6H,14ae2Vg?B&4LSI^?,U6.^5I7A7W5Y#UF:>D5/a;b;.#_#8+R>S
f/)J>JS1E>d-aW>.((=N/K>E4,2E1,gR-g0?QYTWNN6\&#I1^T,Za@^4??GN#+(_
bONW77bT#7>OE3g(2#1Ia_/X,fG27HS?fG,_UaP#W:^[M/(#K#OcP<S([00+PBaS
@f56XQ[UE+/TL+^[3]7-KK>SDIZLBB8UECZK_,.[g5]TNME8OL[ASU136:KH]B)B
@0ZLY<F^C&C>&U[7.JI#1/3HBT-=#4Q5g&D+S5]=Jc[^ab=ITb,B?>bL(.+1C#.Y
Mg9N)&Y3b(U@URKM\b-_TdVe./,eROU[1fAHU=+I2F(3]c;2RgYa/[Z^7Z5eP7-O
NFZN#Z#Lg[=\;b=8)_@_DMDE5S&7M?OVCHP_>bXE^U/>e78EYDWeZN4M)#X)O67g
+4e8D^^WA(BF?/0/THDXH+E<]MGR)cIMNULPX3P_;<g@MG^7/F+</8:5ZMZOGF#3
c[9.LO_]><PNF0;e\#3B3@?8^Fb[O2?JPSa5E;\=FEbV^N^N\Z,/_K9M&,T)S3?)
._U<\H&2G3MgX3C:\e;SAL[F=CdSAZ3@[VQ:XCLCBE8=S@L+bfA^<,XO#fZ@aUeM
E,N77f:UC[+0;A)]bYS;>(E1VRf?A54d(VDH7X&A\gZE=X))Q9Q[W=(HMXc<MLXQ
[F>_Wd?aD-=X(]0T6BMH+)ZE/eZD+WKb:c#8[/&:3]<1#/7\7CR,GLCe&))&/c5f
-bYQ1BD/=^Eab?Y.H+^BB1d[LS-_a\/3>2c,ASNL;S7E[B=_4_#ZD+fLYT-)&VD7
Xb40?7:<YHgSB19:V;)5__.DW.J]5U2>;Y69JSLVV7E)&U=C;T+@?KYN?Y&@cP3J
B[R#BeaY(06.+Q&;dF8fZBFbZ_3+[)20fge+Ic1)a]NEgP=T_P/R2\>eDY8Q\#W0
-)34HC,76Ig+JUVU.5K5.B[8AA(cfP28f98LC4?EQO?-BdVU:-UX0A4X@N>N^D#U
[?9HG+-^#(gZ)3[G,@^Q>4\,.D>#O<)5@PR5d7e;V_I/PfAc5]5YAbI6UU<U@(+[
2eVM#0?+G:e>CSIP=Ta1C:]W?M#Ka]5G@WV03ca#]9P<BZc@><&Rb38TC(\3B)C#
a[]T,17\(R3Wa&,HZ>VcCFIS/JYdMI06bEOQ&\VZ&G5aR2#Of\U.0,#T16E(@=A8
3XJ4\;H.GW56gE1QP2U?E)cdPSH(?U+Xefe)?)]_8+B^CXDNVZ(E=/9U\a;9\I,]
HR4@[@07(T65EK<-U-[\SEVNP,+RX)&&,=2]413^M32dZ&7e?^_4fD<0M1&57;KA
I/14P?d=53;<GW4MDY[=.W.0NTI_<c<C7R344EZ.;F7F/:H#PeVS7&I0ge6C&+:9
M57;VCC<BBg20UGR5^0)6GNADE5J593QMQ9ZKYCbMAgG>(Z-@(2:2A>>=#cZ1UM,
HDH/Y<F?W4O;E@bJZR)IM8^E3]OHE5bG;SP.RUGUSHJW5f&.;93KUZ4Z@H76G>\S
=9)M(74<&ZCUX<I-7?1@&[X)b\>eb1E[-&S0+UF3=fCS[1H=f2V[YZN9a1T5(O3;
IS)f4g>C?cL_LYIKM=gGJ);)DfUCN(JSE=TgCI?A_2R#/f[?-3;DW_=MOKJ\7EK<
+J4a_&S-[7[GR\W#&4#4fL1,8M0b)U:TJ)fD)<_<SSMdVSMQ\e6,97\0#OYdVLQE
bgOa=A2:ZPW(VT5OHV:Y4+N\@37^,Jg+[]DYO;c2SIOPARg#Q#DN:_=(C/H1ZUB9
UJU-J)/b:5[bgc.EC:0V&E;Ug/a(JK\1.cZ63E.A8/>A9_RJ;C_5ED]VY[;GSNRO
g+DG/M.J5D6gVgC[I.XK=IB+E3Da++;bQ6Cb:-ZAZB^P(6U?Tc[_0L.fNP+X?P3(
d80NgOc<@>O8e:I:MM/?MZFGVA1G6^(DDBcYX9S,86QJc7+\H-KNJYW16CYC(5X7
B0MY6:e;2VL3>Q)B>OfHd<]4+Y]LRLU]NF#B[>L:KQ0F0OGPX0FS<Hb<Ef#BDFIR
A7d8dF0.S,-ANe+[PVeEb6SKE3EMc^=V(+7CK8/_TJ^6_>W9]W@a\ed5,(cD?F.:
X4<MVP_4+W1d_/CcPZ)]+3>bJOH195,:<\+#SJ_U)K^Fac==6EU&4DX8I\M@U(D\
W4fcTADgd4)6/-T-4D)D#1P^BW4AGPJ,V-1CRM:SOc4V1G6d,Y9=QE?(agF7DI1T
-EV-&DGZA7I<2XWV;K-1RFZ?HgET,fSKB@2Z97HL4;);]Ea27ISPG67,CT969e=_
f]Z=e<)P8<3JSa_\,eNX^&:3H]H;O9B/?ZE]&4aR@4YW_-95&?73cAMGB8;)@H>A
&200FPFPecdMS8I[W(VZ1?IXP=]2NgV#577C@A/N/_3SEf-HC:d0M[5=ee=+;1Q?
M<UK&ZdKBKe9)F0dfK>78+<=21BRF/3J)0BCY\_+C9P392U06HZ\E:^=WSI#c060
.e8CKX?L2Eaf3+(d7B/84]&KEV,N\U-5eI9a<?@_Rg(#^0=#gM;O<IBN0?8;RDT5
1L5ZZE3[L[)QDL@]Sa5MFZ80R?[@d.+R=[@G5>9+?TS@S\_O.6e:4S>FNIU9:Ae#
=aG5N@+&X9X,V3)#0@G0\\J4,W(@P/3VLZBPKGEF-OdCAQH;L]?CJ5PP(?P6cKTF
Z2d0<W>bDC1eP83TE,(TEBd+74@G03=M)aWbTT8NY&9R5D_LJI=]26F2c([cH?MG
4BA_SfO;)WC+G4[UG\,<d].4ASH6Q@K0e]0].e.P,^EF+\4ETF>KS,_f?WS(L=aP
,D?KW;)A^,C4g^G4]M_YB\\#Y)B13?J#;.^OL+<)?5EYb+2@^:?ZeO3gM3B+)Y5d
b5X(MM60O,CI^D>ZL/GLJ\fQfN+>Ecd>5][ZBTL#TA<7gQN&g5Eg;T+[f0K1GB\M
B=@UVLOQ]?QP?f8??Ee+MF.RVHMKZX/(aX#?WT,0><C:E#G^cGJ5/=4EEY0@M@c/
FC,ZDK:-&L)-YSFLCaJ#O?;>XHL.#]4\gR3d9DIG)9B)T0TB(GG6[/OX=&Ug(bFC
FT_NFLZdbFCa6SgGM7JfJ,G?1^R+d]JJ>+.>=b#<+4@)[3;TJcfa-,3FBNW)R=8I
7<Z:83O^=M?J0MQG#V-+A&#P73_ZF3,IGL/;I4,Da_BR=W4OUOg04f/V)P2g)c_=
DeeTWK)?g@8?R^C5V2DCJBT:7:JC@8.,)\OS)JVW06BMbMd2>1;aD9gN)_H,NJcN
V\Pe9+fWgHb?.$
`endprotected
