`ifdef RTL
    `define CYCLE_TIME 40.0
`endif
`ifdef GATE
    `define CYCLE_TIME 40.0
`endif

`include "../00_TESTBED/pseudo_DRAM.v"
`include "../00_TESTBED/pseudo_SD.v"



module PATTERN
`protected
d>P;g+=2]./+fD\LL0O\5fLL),/]C[SGOfCCSN+@NeJJ2QMeTX9F/)S,dUZT2JX7
_(GGP5&5(#?@2,3RYR:BO_90;MOJ1[IUd@>>D]@([T3]\64(FdCKdJX#d#Ma1O:L
c8T,L?^<=65VWf0gc&K&_<OLYQ:CV2N:<U)gEf8@c/d5aYS?d[3cDY5F__IY#D/Q
UbO8AIc.UWc[M?a8AFE+RIX.RPc\OKE0>de^M)B#LONRP>8H&&=.#,IcA=)DN5f6
d=+IgH[EQfUT1WI_d[.:&(a>P:?Lc?3g1L9LLEf6e)ggS&A(X@>H3QM[P-V<eZPg
?+;;3M)J6<DH#,\1CcYT?OBE]bLU/57?)CAgJg6T>VJKFAPRAVH.3G;0^1X06F2L
GeC(S45H&1-dXU26OIL0+@]V.;CRO=DM/EI8O<U)5,e#Q;<^+:MBH#9V/26LaZ>[
>6H@^D;YT;f/_Ic#4GfX?dV/9b8C^GH5319Tf)FINc,IJaW,#)ON?W[F.+(N?S33
6I82ZV\>V_2eaDd@2ADO^&?>NF+XJ@-#6)Z=.g5+RYe/)OX@d4EFT6Sg<NAG]^K+
c4+3FCc/)U;YLV-N]W2:4J^c:#5cW&HUT=JA[CQ[4f[1A7DJD0B&AdbZ38+]^=2S
71804I7KH6:4,WMBQ=R-;gXH-:].CQ9-PFNDSZ#]:a9O][Ra@@aOO>F^PRgU_7)N
;\X5A6^JDa(B4]X[3d:E]_\I<dK]R&+MZe)bS+:GY&R(:2)R^+_\_0+[B_3+^M0I
(OD<RH+)#XQ_eg#OS\g^WBEV9A@_:)HaY)-HW.UI1c:V/&?0R(\f^K;+T<d\MA@R
0E57<PP\Z5K\X_UQHM<PU&+b9P)2K1WMJXH:M><a)@--QI&_MQ^N-5&^D1,gUQO/
e9S5&?HcH7[M>-_D?4L-4,f03b#:LOWfJf8<dBaM7ZM.X(=bX)1[^W[LZNUa\=,C
0<]Z;;5R?;W>4H5fL9[+S\B@>7>SdS,SA_IdZCAHb9#OQOfK5/L^9]L8[Bb,e#g,
K,+a,X2ZW4B4@_FLF2[O2(5^V+b?9?2AT^D\;FGg<@W2+c^9FBOW,N<&#UU35)Da
NP3T4T41LQKcIAVWV#=[-#M_CS7Q\(MAFKC+5X66?:Ib2HN2RScR^N,AHe2,>#M[
-+2c<;YI2GI_a[X\:>R.->QB;5/WcF-&:Z[0Q&5^bbU<PV.2R44+2\/cMN)f9f>L
LTDAR0)6QJHFE@23;<B/(]CNd-eM:fZIGW_E.8BI^(RG&O/BMYD-R9QA+U:G<+]Z
3caa)LbcY/?6c/C-9L9#3BRQP?ZBO(<UP8B]c1U-GXC[U_5RG)YXb/-AX8#VVU53
SVZA>_WR>BMf<=QcU_BGB::AC]^YHFH-:aYC&EC7&PW#e&I4;59&PdT?:>D[8bSS
X/gaUZN)&I4B:0bS[=c]YHKO#BJ[F(-[f\BB_C6=RPQgY4VI&BI9\bG6QIANg)A3
=4D1,UaC_NQQEWGff@XI1eU,H+bHR2UQNYBL0P23@9^+1-5e>_,>)PC+G7#_)BB-
/&3L@F9J&Q7\NZ?ANR>7D)d:Y+9dLUF^=K\RVe^bVEb/#7O\2AHUa#<7_J[bgZ_/
CG)K3VV+PVBJG:(AX#KcKN;+Md(b8eN0P)d#0)/HG>bC>A#\Ab#/]OX.M0(Ub:c=
Z39a.<P&<61M^Q[FX.<M3+d/_1&/W&U9<XUA=ZAbC^J4L2C,UU?-fdgMW2:g8R)O
_?PM:d0]-\^@[&GcFf=-G0S@]cY4Gab-Lg\7V3g75?K^^_(,<K)S4J?NQPBb07KS
\7AGA?PR#fe)M0PYH5K6d1T.bY&110V1HW6SXX:f))./Q:ZTSS_/0XDV6Xaga>TR
?E5O]X_LPN=SfB3B6W;d\Q0(6:#Ga9cF7P:PZPLJRC&@X]X:DS#+A0<2Q_#JPHS0
MT#e7=TObA^:YU.&@M#R\&:X1D^@13VY++OA-?UgMJ0=UN;EFC^?XHdFG&89^J#O
;X(eT0=?0)dI6D>OTJPGN&.1#784(f84.Q)ZHcD:,@(BM(\)<\N79-/&SdEO\(OS
/+4d\M)[[W=(G[MJA\YDd>;Vgg@CLL7AKb>\=WH;)C-TQ?e\Z(0>I5Pcd:M8L23Z
/SUO(&]68]9<QG7\9_7I[V&RAK42ASE-NfJ^T\Lg,Zg;bNP828P[=_a62R)K[+)#
&1Pcfg_>N55d_;b+Q::N\:H)>.)Q6MHCJX#UG8,0K4GOF_aQC->J?U-d8<4fc\I;
?OPTCf_MS#;,R:Z6CHgaSK]K:_^1.);_[(Y?>(\G7]6VWGV\)?_3(C-egaa3.T(f
6<e[3@M/[/,C8RTUZ?BZ1?.=Q71.5<3BC,>6P#N]?2c>3\0ULc?Z)B[M0/(6dgD;
BbX:R81UVVE/4.8+JZ>=?B<8<EG#Ka&bCGX<XGLb1YcM.+egI2f(=0c0+PU-#=NR
#VVV(Sf9e-^d4+6398Ue^]M8J[/8(b4=;P\W<6W?-Q&-.Y>8ad3O#3;6Gb#D:W6G
)R7?I?</<fF24b0VBGLLK(@=2K-Vb>g_<6YM:eN5.dB2Y.bXLJNf,VTd6G7H/\Fc
K28Fb37ZbF1Q?&VbPTE6?0I46T[KY;_565D:Q#g\0IDJ9W?,e=)5G8\N_<;N,NWd
Y+JN=fDX[-ReWP9\3@f2bbdZ;-PSY:f2_;A]?\:>L_Gg8:SeW.EVVY-1c;Ug^f&\
K(&F,YB.,I&gUbOI@S11\5b4?=JKY-(?PYe74&?[=9(E6L#648PVO)?;/L/KX<S:
).&Vb7BZ;9Y6+.GcWF#@9eE>\,2X4L1(eWAbO@e^/+&N<3AE4;76O[32LVg8WFA4
)/=SH4;fQ0V.f1V@VN,PV4<-2d\c\9I1Yff2+b<BR_eU1+?ZS7Y)7eSVd#;eJ9gM
_2Cdd[GRGHDKW;F=5WNTc0/^6<(HCC[1R>Fb-.KB[a_6(C?JHJK\e^(&FMa>5cJI
8H/(eKJ)>Y.CCR_:eE9gFW-8B1fAL2Ce@C=ePTZ+3H4R)4(7SaY+9X/)0>).B]5^
>cac+C5A0gORAB?51(\EK]:20XTD+.,-+-(5@RS4eG0)_Efa+b9@5]GZWWN7S</@
/VNdHU_RZMb9YM=QXL-),_.W?&C&BHH)aAFGLSRP,9#NEg13,POR_@d#aPa(6AW,
4LK(J16g6S1^N&0_MdH6E+.b3a68@J([G9T;2#>I+;T?dBSVI15ZP_dZg0Te@.A(
J_-FNa+;VPg52]7Xe+)+6bA3F4aPRCeaD&U?H##C/,RT6A+_+[KM^g:bY4BN#ZPX
N6XV8X?Ybc4HNG(B[OE+Y5EF+eBS9V)C,5U=d6V(S64f=\S:EZ76Cc^Hef4bF[\a
Z]V.O69.F,/2U4R+7eF=aLS:04g,?8]:D=E&#8CN9@J,Fb.A:+R>fc&343c+/UbP
V9fEUW0[D//O4faUe-a9G)5,>E@V157F<+;S_e6-3@3EbfBeNW?O^d6EaQ>VGJ]W
@V13/=?P+W9H9=1W9.FXZR?WCPH]^M(;7M3+2KBW=dfdI5f/)/QTc4I5@,C^JSL0
GMDUKT(R9<gX9f\/LBC7\9L:(dMTVT#]Qc_M).&Y<(K3O./TbI_UY,;dZ#Q6GA;W
U#I/c+d3^;4.;(UaVdf^N87<HP0L[V.N.&QUa;XGVX/(1MP^RS,HD9=GLa-F;9\V
BE4L\XI,^68))8QAPL.E.L#fVB7fKIfaIQSP3RV3SK-fQUXK@CV1M?CVA8Y?9agM
T-I;)DXD7N(?25HHBdF3:/BPQ_IPG.D1IS=E6gPfBFW^OJ25OBPGR2P5\<04/P^?
C]0D&SdCSV=cIC[A;X^1g2B=>2A2Fa#T,YYO/cbFKcBTHJ4^L:2=+D.O@-61a=2>
R\dA8Z??^^:fHMcgJ-:SSf46#N-G@H3KE;CZ8cc_#L/_Ae&_1HUA4#N-T\+.GW+I
WGe2?.S8(G,X\;=f2#NES>C]dJT4ReL7FHM7<QCOJ=:?K0.4(HZQNLY5P3[cc_SI
?2(0(1/CO^:4&>]ZLYa?WNA2^b];L9EQBePEC3:@b(\>CJNW/Ieca?2/eHCGRF&T
:;,53FGZVeG6Z:&T).KI&RAgW8;0,C18]FDVVZL2_C0P0;dG^+=fBV#g_SD/M08G
gB2<4Ha;IC=U>+NF3e>K6(M_>-NO+fB/RY+<d1ZT0Sd,ENW2A)>BaUR<&/6>L)4H
VgXXT^[PEXIW=HH+5=@\\[cfD?:\dGN6XJI<M7<,_KV]IS9:_ecd4:=Oc7BH4b?.
>Bc[<7#A>;?Y/Nea==NEGd5>(^0.>M?RV6P3NEGI;:R.b,O:b^XEE+?VdR^UJ>7c
\=:O_cQ60d#SL[C:.7=9]MDHVRC]P;VVL=98>a=T?S]L4=aCGK.T=P<7M@WEgD)Z
f?3,[3=bG93]ONf464#/Ob7?gOQ+cI?5-UF->]/\@1DY]NCe19J/WG/=U2^(_>+L
G=W=QAf>CIbTMGcEgMR\[;L;=;X)_CUU2_+S/E0837@H^KMS>eDe3d?X0PDMeU8H
,1SFg?_@e+aSa=(#WPO<.\f.1b+L_CbIV?7LX\#,/g<;KR.A@H(a6,KD9/E.g,2;
W<_.Z+@&TXU>&SNGC7fC?9=WEV^56.9e(62bb(gKK0A:H9f_6.f__H7T)O1043^e
WfRK=4INWggNW+4_;/P[[]N=L#<ZF?RL(FV:c;MIF6eA,P:0\HE@LV6-[b;dHgVf
E-+VD0E+\R[HXXN_8dV)U/]HGYG=RM6^9S<cJ/E@4X]@9>=RAEe<5^\>KCXdRNZ6
:fVM1B-,d;7#ZF?1R@XTL2;Qf7[=?CJA@@aY:<Q<^PF/<W/C8g^]&;e2E9g)OA21
F2FEbOTF03GcLeIc-12=MO92MIaHJNeT2A1PI/(9GRE@T<]+M(_:JSe5SCZ8g7<F
C@BU1d#.6PIS#WR,UMV[<L2_X>3I?/c#5,M:SSOI-F:<HL9dO2?Cf<c:Tc@KGZRA
QgIPU6U=>J,G0<b?d3]\@UKEU,0)cAEZ2Q2.(J,SET6+g]#7)McK-dHN+\PdcgP4
N_J5^HW#QSeAUT]Hf:dU0:@?baNUNM#V9ZEAICJFE3,)#HR1##K#WaJ>E#DTZ10V
2Xe0Kc<f[&<)fe6ED)SVGVY22<DZSP\&gbP55@]ccTZbRC7eVVg?-5?8QL/V]Y8f
;KY#S;&bI6Q:&E7FaV4Z[1D6f^K9.<[ROLPYfVMGBbYP[&H@b=7HSG@POd<SZIZ5
:W3\QE=2@-W5_B&)P?<4fEgTUM/0U+NVc.4/@V[)\XD_\d&[HR(4CONWLc,J1?8M
8f[AGOWYY2fZQD#7\.1R&9X[IIU5fHLB9Y+24WD7^gQ)ARO.X\d2KOE)7,X7_LGK
X4F/V7=8]DZJ6aLI4(PK.=M\_Gd?P-8+(AEdcDE\)U-DbHLB]Td[&DK)5F8+1f<,
]R^]a^9Cf53B2#TUY_gfF2#.>6KO=_B-)11[^fdE:eH&:#4F)QTZHCWc[Ad[c)P]
>1BA/>b@S=#GJ])0NC,&P.;11a9+QTc^cgHgE#FZFcSMc7:gDPM<,PPeA@.T]2]G
<]eUH7b.ZQS2Gb0RT&R-)[;a#eEc,#O(J]Q.5<=Had3BOa5(#O-)722YZ;1V&-/]
_g^DMD3Y_.ebRDUF<);^A9;Bc==<K<WJ>:BT09cM#fA(69HFYAYPge,33:R]LHK[
W+bM/d+&]UaV.gA5cAL]eR60(2PCCNB=7#)Q>6@f4E8.)GJaT2ZbZ.>99#&>?TC0
?M.:fHHP#L,DMSU>6/2J>D[<M9MG7fe@VT_;K<W:8:<)=^Zb.2?WQJCg_ADZTE[(
@D2:@E;QEQSc4g8:MW:PJL[[QH-GIGU[=1g2OM?P2?TRQN.G_T3)-aCOaTRdU+2,
:.G4AAd5@OWd\</d4#WaMWMccg,SRV(=IG/EE:AGE9^Jg[69V/XZL_[WJ\V+XN)g
;bY\P11F[.3F7OU=AN-<6=[]]^^G3;6>71[EA;MNO(JO9@fX4BKV(/Y0Q/(2JR,\
/,X_W=]4\EZ46SQ3]]E@<XN6PR.2gO]])aLU00gaAK^X?WY2TNC@)1J,FQR7^PDL
9/5R#,b:eb4O3SK1K4[/(70EA&->LZIIa@74G6B.VgU\XJG?Gf:FQJ+3d3G<O^O\
S=-X38f0\_._.CD_B-KF_;;Y>BfWCY0S[XX4B869<d/g]MNC]5b^TM:UOSEZJE/K
2P?_^BJIfTG3^KdeB7RI:</XC55Q?;:a3AJI23Kd83cJM96FQE87O@;(,bYNeO+d
<FR5,0f.D6gE?.N-Xf>?P)6dU(e7LEB8W1==W(NFD;_^YAN@=]TbA9MAe^5Ke3H\
J5S[3HTLcQ9A\#Sb#-&261X.E[ZLA;INd,#43?DGTH-JNP3E:d9Y7Q,KR;]SC]\,
\S6TF653NIIf7ZD/e<_2cb(FQ.A?:\_5^,A(&<c)8QR[_]/#FeYVaC/<X^8W@F2)
UU.0?,0Q.4eOMK?,J]ICU31b_c9=PcZ502L@=].Q>&B<_[>LF=g3fObE\<9d2W(/
K<L3eO=3@Jd]J>T6]gZg]6dQO[b1:SHIFM],2Pb?c;V5c0E=M=^(XK<f21\+fD,-
c(OD9B\70=@-949gW1IK.:@RIfc_Q&.G@YR2_f.8F?=CYKT;<8RD;;_XSbK4Rf>^
#&3Kea/bJM-/,-,RcKBf-B>_ZNTT(e-3#>PBg5.LZH+OTIKXd&Vb1)9;fR/&f-)<
,cE&(G]O>4>6e,4I=d2(a^He:_bRfY5aRfde/S2I@^bZg2REcVb+9NGP=?[5)9S[
=KUAW]J#SbTB8@[V);PROQ2\M68Bf:_BWGHVbXCSJN+SI=C4OOVc<g:IK]bEQ8JA
5J(NZS;,^_PTHV7@>eQ19?5_aG.AE?WT9\,VcDBgUgQ(dP25IBELZ^>]LOI)TBK8
V^XVG1GOcSSLYY]?V#4CNGR4JW#W8S]#+B6;7/RE4F[@Z(UNfF7Pd_d#R0]bJ:JA
?[J(aRF8N\QgOgI:A<=9;:dDf(/3;\;&O#-.\DFd=[T@KS+LX_&U60=UPN9H^fN.
1,UB<9T/aJLJM>gE0I>I=G^O:S-[f+g>EI3JE0:TL@:[FRSAFC7Ueg;:NUD3b^IU
<WaYNT1IUIR8cW1[UBe:DWAUH-Ha:R:IS36)-3EQ/.@EX/N/167;OO(YgNb=6J+1
RHO(EYEMBe+_4H29.f-6X(PSZ-Y@g:,(:KL82[-c)c0L\A3EZ(a7g1(4;E3?BZ[Z
N+K:J5dYF@LA788Za1WXYR#>?KUOaaN\<2Z5R;<IY=:OK:G]1+>Gg,=_e1XL)<@H
X6RX@eLBcSJ8^?Qf[DL1dR(1L#.<c\g+OaE73)?5JfQ+(SH8;^Vd3LUK@O7VQ_PC
HPLXPE\SKG^;Ne7d?Yg\G#WB_73#E)K+UZ)P=P?9OZ5PX&,PQ-V;g]#\7DCW^F_H
BP\G-U]9+PXCcX5/RF(;Y(4gX[U5G)5,_S]4>/]..YJ?K58R&_#TAF8I1:fUcU>Q
OLf=7YGc]+#:,^EEN3P8E=4O^e+_HZeUcMg)D6E@6Z23]6NDUSUc(AIWSb_6^CC9
g,HKJfdPC8e[8d+SI=3+?LOM7I[V,QT/gO7Y-R?aE[=WRUA,,X/T>K2AW^Z](@)E
/BWJ/<E=#?e?4?>Y1O?Y@7?=M:ID+5RZX:R[<8d+;_-;b8HV9/9@?K3[MR[HMJ@X
+9O46SdaE)\7\VCV&V1K@Y<McP5b_YbWDUB&9;^XH1G1CY<Ofd/EW(>?b>3#>;8D
>EI=I>gea16df?#5+A?eM<<CN4+Q<\^.>,U(&-+S)<JIb2_:MNNS4#g9W:RQ-gF.
2S?+)RNT@),^ge&6>_<#UPU,.&(FR967UYV@:.4@&76Y-#fKU??bHC33U#YVYOVM
)5G2M1aJO(P.(JS7PXg=8?XO?HM4EB@WH0V2a8;N8I)C/N,F8;L<@TfcQ#M&KGA7
\8QfDfQfYVdP^CDYD8+5RGXOGV=.Q=_/=^1e?9=WY;g;Fd)b1HaX2O,1R?=4SW-6
4C^N>-,P1H)]OIF7.e&M+XFaK,N_bKYQV(?NWfHKSF:YAcbLYO>588A?(38113[=
43D]32SJY(<[\KEP:=N&()&KBH=^)E_-5f:L_?ZL#P)](CLEEYK/)+][F_\:;>=N
G@S:>M5R,K?fee_;/eJ9X7VEP#KMc)M?8BHA4@;]/SXd1TLA1LbL^]K@9S=QX&[>
0794-JP^e3:Ra^\a(c7geKb,fWc=HWD6?DN-P^><bKJ7NQ654GLd(gEJCPQF[R/f
H=_N#;8Z)K3AR&;ROMID;)e=U6Y2.BR3RDTd]#:=7TY2BCH2BLfGOc,gDg1<GdJ:
ZGgGRO(\((>5KB07H9)RN7IdWKW3b8dYdBC6d2KPI<3dYe(J^DP-OG_ZS3S-/\OB
GD\8MLdg/LCSY4F^QSR4N;UV1H?F)Y)cQL4c>(K-<@3>E,7GWf6/2cQ>a\^-[JP=
DTN_\B[GcRJ:&Ja5NYOET;d&4#XMe;=P;DPa92A=Gfc_8U78O1TQT&+=WZM2e+U[
(D3E?_B3\ACdH2IG-Z]Y+YA\:8cX299Xg2K9,WdH)]W-C^F7ZEf@<X29^.L_TU.f
c]PY0H?96S3?67^Ae11SK(S_/5f_M+^ePe+9S^0LEK&AY0;Z(0URY9D/NeS6E-cc
==_8fe\WDFWJ_d:D9LaF?F(9e<\K4@D3V,R>YgcTS0KAUCf.&@a\]#PQAaU</<2O
TGLfA^UF<@Y-;8AUg0Ybb=5^3-^C2;6fdG0[c1[@E\ESLKXH#L+EQgNI>MgTRf#L
83,#JJ+YRMRP7#S(-e-SF;]U[<WC>J9T&@RO#g_WXQS>6(3Oc0Z/@3FI/<UXEW)3
4bdQ>O_Y&DPT8fFZ3.^-dDQ\R-fAdJCY#N99Mc>Y-DJH<07_XTCQZQ^abULf&b4I
-a/SdPODD^??D_H.:V9>P-cTD\B^JWF=GcK>G:0&f:G9WZF,g#N]U3/+,f,E6D-(
HBSOg;V&0H-UMEKf2DRAYT7T.F>=<gOgae)ZXK8TVPVUH<KbDfDX9M\H[N4;7g9H
d6Ye_.L8V])YOB9D?>#3ON5,[OJ-(<S35gX\]K^N;19H<c00?g([Lb1R;<+5fG_)
6#5@>2-GW]2AZ.Bd?]b&eWMA).=K/]7(WeD[I67ZQO</]JN;V/c55HAe:)K4_4GW
#A^7V?JL#EB,J^10(<@Me+RMO0+K:#?F-gX^f.F>=e4c)D&<\LdYFJDU.9>d(7>,
/16&U?cAAO(0\I<U[)UUg1,(g-Q&5]NGNg.K^9L^[LCc6B6Zde7)\f2AV+,J/+3E
7G++4LXf50,?V+AM2KNPMX^1#-/<(NAcY[9X?51@JG#B8X\B+f_\,:V-SFT_e_^R
H;2YUf>)&#Nc7c+)Q9ON^YLc>NN#[(_2?=KKBVZ4I1.;W<\FC-2?DQD8J)4Y^KNP
-4?HfVV8V(0N3Tf^#_&P>D,RWRIDN#_Y@C0IKQX04LUagVQA)&1;-BgO?7d-Q7eb
]c+Z=cMIaX0-Z\Q?AVS26R8EO)X4_eI.F-#e^4R[7HV0.\.>c3a/63[W]\bc[KXa
gC&C2e<^eAee9>TKIH>fO=&0RMTbQ#g3&^-(MVN/A(aA0X[+&:8g](cR<_R5+cD3
HAeZ;M^T3YXb8(M6dY7GB_fb;35KSY00EZ0-X;M)5Pc)SB1A1D&ZaN3d4?^7X7HY
]VWg#H06TH&OAF@RgDfPR&]7&3.6<V4=6+LHJ[P-0[MAUMUAf6\V+7SeK:&-TT.O
O-QHAR_YJ3ff9&LFb0U\5Q;+/-S_OBL8OP/Z+ZP?0d:;-cHLW<L;&WH\LII42P27
R?9Y;0F8=_FY_EdOZE4W9CL.A9R62>.4_O9IbO[?A<E>gUbd\H3RG4YOWKCEJ&BN
4MTAd<)2X</A#[MCfg);]AAH_\Q^YHRc,b6G8L&>f)0=PW&Z0UbC5(N#IO:PU)K/
?G6APUg=J/2^+86)[?^;=MIN:M1T>>R@8F;#1ZDg1J1[FEe[d96)1e03bY_>d_<c
Z,BaYHH^KJ9/X\#5A#U6.f3E12\(8UKBT;cTfLc0-D8_Y+29-X=GC#]0a-Z4_+NQ
XVT]2H,Nfba]:MTf.+2G(_AJ8AP,^_<8AZPKVd-fY:-X+,ETaS3^IK-@U:BD9_ON
(GZ11(a4cZT^Kb=F[5F,3&e?gHB=2CSGM8HeCQ6#S[M.B)DSS&\14a.fgGgbTfd=
1XAJ&9CVS(J8)I9SbGSZBVW1;fRf/5L;=bM>7SfQ\39:Y7RBMP;=8\<;b44.P3V,
>GF:-+MFNWSM[3gZ0c:DIF\)3C>NAN.(JKT,(/[[Z8:gd3S:#X=3CVDX.5G(g#B@
f8Q(GLPB3aRLW+KRVf9N->7eNMSAP3<aM_RX#)MU@^4Y4E+Hg+U](.3&EB#DC[7f
MH(FLEg::+g3]fTVBM\b_B;:W@^4;916DWR#\ZSF7JDc4O<):d<7CZScKM,^:>O+
78#X=YB=/C.H9P]4CDeV5HA)E<23ITAR:]d2_WS)4C08F95Nef1d6eaf]CfMLfdT
AXMV<:bALdB<D<J7Q7;?6CCGb06M_M8M&6SW@5<RC5SCO13SL77eB&E<+1?O(/g?
<eDVLW@VcH-L)f1=?0Uf4@:,GFF=E4=aAIg[1dd+2gb:X1M4(Y;?05fN#)WO+7;@
DGY[6(CO,4EH2DA;5)UZ20]Qb-4=5a6a[1Q@S4[OS&^T7#TgRZE\3J7H[)3a^a+F
G1A)>]3cLR]YIURMD+PHKN[00II[Y]XI_f_-]Y1CK3?a5OLR?eS\35Z,;&O,-W65
T;N?6a.>__/,4PB_LA2@]L+?KH@gH]CH-DS.OT(/;R-O+C:cc4+/M(,B;I2=A@7,
#LK1Z=Z+>cMdef:aXOfDMgZ-3,d32QWIMf0[:K1_UHMIM>eY2L[B#=[IdeT5UO\8
O^ML(=BYVPQAf]W#959HK:=_//9^NCCE+X6?4=cMHHNID))M4@&HCI+X;d#5)>H0
]/;>;_Z[,eDK1PS)Gg1.#HaW/dT46K1c:PWP2WaSdg\2@8;.9P/4^F478[&SAV&_
gbNNQBHT4^)Ie7=X;_cU2YCaSL&>L^;&egGCPX9VD9aXO5S4W9N>/f7U<2.\&W;<
\-b_<K((;2O/OS,1dY,)\ZRfUc.I;UQ4AL8[)4Z[VULef_WFMc,^7HMI)Z(UG8YN
N:<c2c^?d?:4Q2@P1QKY4ZY+=g_OSaF&U#H3W5W)EeeK:21MGdT^B0YQ6Z@G:]Z^
IY5XJ\8dS\,6)DT(d3/e^2\]AJ+CeI=aWP:+((2(AYbEF512FbYM9U[,=)W-:0.f
35b)N,fQc2T<^B17K<aQ#d0#W1gMB#a#KHI>VG,TN?SZ<A.//T1UO53]YWcgYbd(
07>_BLLb()^W/g]_7@UHXgK>RUY&FZYO<RfL9L>3\U:6#<Tf0_aJ<G2#07]#QCJK
8U4=#=-aWfUMB4R>026a)#D8<#dJSFdTWZ^#TYKfeg]JFLWec@S(\OUD=G035-_a
-0FQ_(1WPNg;b>A=FMP(.=:<(20XE5Z:FO@E\J^gIK+I->cc[:ed7C)GBE>bQ15F
AN3B;1D)?5?8IYY0\))8#[PSGJaND]VJO.&(WR_=A__eEV;<19&7dMd#<gKD>;GK
R3C])<5X@bHQH_P^-.?,3?>[c5EWHK-(2&)>,9cF2@A(&]EXNg]@[8feRXK+c)9[
M6X^4eQJ]J0)AVXIAX+C-WZJ6\&Rb;&P#Z&(1fe?N<Rd?<)Ef4V\(9QeAKIMI3Y,
QH(b/-=7,]5<L1c7+Ua2@[3>25Y4.FC3NEYTFNe9.5+2>X.Sb]cET_MRE8+,\aAN
L,6ZeMO;Nb<:e^ASUP1d[WY\K<O<.GUE,>DXgHb;cE<QFV_6UB-]9WR97LR5VbSG
F?c0UK-8daK+S@]YMb3;Ea-&B.OTQHP]]QbR/c[UPf;1Jgb-+TeSA<F]Y3G14JYP
,&FAJV87JE_c9#CVQ<cY:@4W(gW0N/(V>U5,,W=WA,Y)O+g\G(;&UeU3b\0g5/,8
LEX;X-5FSQ18Z9QS=;RcSO>ccS]7A(AJQ^2WYRFV@.fWDZ/]17:]&32UWWMGWULb
MIP@fa,b.PX5,U-:1Mgaf_Wg/6USG[&,c8_WX\<&7gYM3LGE7YZK8NA,EE./+aZR
fFJca;Mg\_R3EcY&J5F3;/GBN<eE^&@cSI/CP6=UJWG(KTdg2A;eaU8A<>=1N;#G
6d(e\dgEIDUg30?fP1\Ef@=]dJ+PTTL0.&#:/<\>;^;WIV_SgSc\4Ac_-IYSJ2CK
\[<-QM>>6UMd54_aZaaI@]?.U-b(<>@N#J5H]d5]+>9RaD;8#==bH^J#HPY146=,
F7RWB-2XaYU@/MQ,7e.<)M6U/JK;F6U37TG+)D8G/I<>MBX^-U.?a#2D7^RR=)+R
)U^Q_\7bQ,Gf1:.>#JK#9.bC_JeN2D\M21GN3/6..ULE]8(8XOBc4_3X#Y-bg>0.
FAUM2;=MbX-]LB2cNeRSHBbAK6^E.>8@\#)+@A;S/3I;N^TQ-@D5[<Yd17g#+c2B
_)^7HO8:LKZBUA1.ZNH6&X+1(e>K<GFW#/R=(I3\I6.;_CCG)_TE9=M@#Aa2<A_+
Xf@P(F@S3^g#FDH/):9IP#O-T&6VX5]W^GbC6)3VEX3Q,2)R6:D#<M;LQ&c^O(F9
-6P_JI;[ZEN5FVX\GPE_JE5^X[5C_IUdO.(45AVa18S,SVN:1_,:0(X<_N<113b:
ZU5L4d_D6Ya_3DJ:9:M+5f)+bPE-.Wc5-FWbecQ56P3M0P9]^77fd\2E&f\40[>#
AD;I69-e/Ge1]+=;P]#BLf9OXOdZX<?38f;9(;L&WN]&;3IU1;4FG<#LOE)+X>.8
=b0:7GC;O]6\b2(TbT,3UL3FICRIaMB69cK=C#4#NJ??/4&\EeM.TK^^M?7:C)f5
^86c:3HDF7]7RW)/4aPJCYb=)F#GT?E:-H2_gLY7P(/^Bc)/:Y\-[L\Xb]d5Q<YL
d(KXKYcB\NE5K8MTF/dGP>>4-?TEP0T-b+/e9M;0bE:Y0AgFE>);BPTG:Qg=U&&N
63S9/(C/L0:SFQPLaNdYY2>XR)c@E]d[=Tf+_9.VOH1N)28PTGd;/^7_8JN5aK,R
TB#T8eE(9&geN_X)63<Ha6C6:BdgRFE;eF0P>.()/L8f+6RCNbb5FbN9d,X1U4RB
J1&QL904G/6H<b1]XGS/9>J:TU#C[S\d0V0VZ:^0f<&N=EIZ?).KZZbS-AYc+1dC
B,I_S:bTcEc]6M1.JOHB1;LdP>\AHZAdGI]I59)8?;E0#6JGKI42+=IP-Eg#4V[K
d=H&53\[PJS]L0ZV2+.&M.CMgfe;14f2@55H^36&CSJ&B2F&7,5Ug54f)(;M,^\b
.\a:d@_E]aA.X2Q7+33A[4S0NJ]5RS;bMbWF^Q\<)1U:5&V2C/Q@cL);[_557Cd6
MX<Jg#);(]0ACaP>@4CW618Id)fG?\35C#4.]2dCA_W\9cD@)6VT-DJ2_.g1V.R1
]E5[ZRIYZ3UL_a)JYC3aNf7T/Y&[c;Ec_VR8D,fF]>)YDN[R/=:CH7#IB\)dA[I&
AD>BTGTd\eG+=WR07#K&K6D[U4W..GN[IX6ffA7CGMV12W#S&X(fe+f3/bP=dCN.
85J4b#3cY<@3R>Z8_ae^D-VBS\Y;#RGG6B1ZdL#cOg[_Lc[Z=(0e?:1+3DPNM@1B
ZC?+e^C][X9_N_WeK)N;YUVS+8W3J>fdP5&I2[\7G)W,c3La#-+cG8A0Je:JR6ZH
;4cb/6[^dOaO4BRC2<CQQ,EUP\S9?EZP^S)b2:D>/>b\^6]L.c2fUA/<XfVK>c]+
&CKM6MF29X1.d9<bJ7XSQI:=UZ_4T.&GA@&\OE.)S@N:I]V#EZb<CF51Y5+^N&F.
_ZILIUSDZF_K?;&3fbL(2-E2/GW;F+RAW\]T=.TC=QSOJ@V.)Q.[,2F=e9U,)Y;Y
5f=RO[7YU=5)7U-QZ-Y-Cc6eFE7)9=D;.0KBQ[g7L+&I;<<7JRSC\0F=J$
`endprotected
endmodule